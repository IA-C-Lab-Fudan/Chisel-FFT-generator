module Hanning(
  input         clock,
  input         reset,
  output        io_signal_ready,
  input         io_signal_valid,
  input  [31:0] io_signal_bits_value,
  output        io_cosines_ready,
  input         io_cosines_valid,
  input  [31:0] io_cosines_bits_value,
  input         io_HanningSignal_ready,
  output        io_HanningSignal_valid,
  output [31:0] io_HanningSignal_bits_value
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cosinesbank_value [0:719]; // @[Hanning.scala 22:28]
  wire [31:0] cosinesbank_value__T_32_data; // @[Hanning.scala 22:28]
  wire [9:0] cosinesbank_value__T_32_addr; // @[Hanning.scala 22:28]
  wire [31:0] cosinesbank_value__T_4_data; // @[Hanning.scala 22:28]
  wire [9:0] cosinesbank_value__T_4_addr; // @[Hanning.scala 22:28]
  wire  cosinesbank_value__T_4_mask; // @[Hanning.scala 22:28]
  wire  cosinesbank_value__T_4_en; // @[Hanning.scala 22:28]
  reg [31:0] cosinesbank_wcnt; // @[Hanning.scala 23:33]
  reg [31:0] cosinesbank_rcnt; // @[Hanning.scala 24:33]
  wire  _T = io_cosines_valid & io_cosines_ready; // @[Hanning.scala 25:25]
  wire [31:0] _T_2 = cosinesbank_wcnt + 32'h1; // @[Hanning.scala 26:42]
  wire  _T_5 = cosinesbank_wcnt < 32'h2d0; // @[Hanning.scala 29:61]
  reg [1:0] state; // @[Hanning.scala 33:22]
  wire  _T_7 = state == 2'h0; // @[Hanning.scala 35:14]
  wire  _T_8 = io_signal_valid & io_signal_ready; // @[Hanning.scala 36:26]
  wire  _T_9 = cosinesbank_rcnt < 32'h140; // @[Hanning.scala 36:64]
  wire  _T_10 = _T_8 & _T_9; // @[Hanning.scala 36:45]
  wire  _T_12 = cosinesbank_rcnt < 32'h200; // @[Hanning.scala 38:70]
  wire  _T_13 = _T_8 & _T_12; // @[Hanning.scala 38:51]
  wire  _T_14 = state == 2'h1; // @[Hanning.scala 41:20]
  wire  _T_21 = state == 2'h2; // @[Hanning.scala 49:20]
  wire  _T_22 = io_HanningSignal_ready & io_HanningSignal_valid; // @[Hanning.scala 50:35]
  wire  _T_24 = _T_22 & _T_12; // @[Hanning.scala 50:61]
  reg [31:0] hanning_signal_value; // @[Hanning.scala 57:27]
  wire  _T_26 = io_HanningSignal_ready & io_signal_valid; // @[Hanning.scala 62:47]
  wire  _T_27 = cosinesbank_rcnt == 32'h201; // @[Hanning.scala 64:27]
  wire [31:0] _T_30 = cosinesbank_rcnt + 32'h1; // @[Hanning.scala 66:42]
  wire [63:0] _T_33 = $signed(io_signal_bits_value) * $signed(cosinesbank_value__T_32_data); // @[Hanning.scala 67:50]
  wire [31:0] _GEN_16 = _T_21 ? $signed(32'sh0) : $signed(hanning_signal_value); // @[Hanning.scala 70:37]
  wire  _GEN_17 = _T_21 ? 1'h0 : 1'h1; // @[Hanning.scala 70:37]
  wire [47:0] _GEN_33 = {$signed(_GEN_16), 16'h0}; // @[Hanning.scala 65:32]
  wire [63:0] _GEN_23 = _T_14 ? $signed(_T_33) : $signed({{16{_GEN_33[47]}},_GEN_33}); // @[Hanning.scala 65:32]
  wire  _GEN_24 = _T_14 ? io_HanningSignal_ready : _GEN_17; // @[Hanning.scala 65:32]
  wire  _GEN_25 = _T_14 | _T_21; // @[Hanning.scala 65:32]
  wire [47:0] _GEN_34 = {$signed(hanning_signal_value), 16'h0}; // @[Hanning.scala 61:25]
  wire [63:0] _GEN_32 = _T_7 ? $signed({{16{_GEN_34[47]}},_GEN_34}) : $signed(_GEN_23); // @[Hanning.scala 61:25]
  wire [47:0] _GEN_35 = _GEN_32[63:16]; // @[Hanning.scala 67:26 Hanning.scala 72:26]
  assign cosinesbank_value__T_32_addr = cosinesbank_rcnt[9:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign cosinesbank_value__T_32_data = cosinesbank_value[cosinesbank_value__T_32_addr]; // @[Hanning.scala 22:28]
  `else
  assign cosinesbank_value__T_32_data = cosinesbank_value__T_32_addr >= 10'h2d0 ? _RAND_1[31:0] : cosinesbank_value[cosinesbank_value__T_32_addr]; // @[Hanning.scala 22:28]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign cosinesbank_value__T_4_data = io_cosines_bits_value;
  assign cosinesbank_value__T_4_addr = cosinesbank_wcnt[9:0];
  assign cosinesbank_value__T_4_mask = 1'h1;
  assign cosinesbank_value__T_4_en = io_cosines_valid & io_cosines_ready;
  assign io_signal_ready = _T_7 ? _T_26 : _GEN_24; // @[Hanning.scala 62:21 Hanning.scala 68:21 Hanning.scala 73:21 Hanning.scala 76:21]
  assign io_cosines_ready = io_cosines_valid & _T_5; // @[Hanning.scala 29:20]
  assign io_HanningSignal_valid = _T_7 ? 1'h0 : _GEN_25; // @[Hanning.scala 63:28 Hanning.scala 69:28 Hanning.scala 74:28 Hanning.scala 77:28]
  assign io_HanningSignal_bits_value = hanning_signal_value; // @[Hanning.scala 59:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 720; initvar = initvar+1)
    cosinesbank_value[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cosinesbank_wcnt = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cosinesbank_rcnt = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  hanning_signal_value = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(cosinesbank_value__T_4_en & cosinesbank_value__T_4_mask) begin
      cosinesbank_value[cosinesbank_value__T_4_addr] <= cosinesbank_value__T_4_data; // @[Hanning.scala 22:28]
    end
    if (reset) begin
      cosinesbank_wcnt <= 32'h0;
    end else if (_T) begin
      cosinesbank_wcnt <= _T_2;
    end
    if (reset) begin
      cosinesbank_rcnt <= 32'h0;
    end else if (_T_7) begin
      if (_T_27) begin
        cosinesbank_rcnt <= 32'h0;
      end
    end else if (_T_14) begin
      cosinesbank_rcnt <= _T_30;
    end else if (_T_21) begin
      cosinesbank_rcnt <= _T_30;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_7) begin
      if (_T_10) begin
        state <= 2'h1;
      end else if (_T_13) begin
        state <= 2'h2;
      end
    end else if (_T_14) begin
      if (_T_10) begin
        state <= 2'h1;
      end else if (_T_13) begin
        state <= 2'h2;
      end else begin
        state <= 2'h0;
      end
    end else if (_T_21) begin
      if (_T_24) begin
        state <= 2'h2;
      end else begin
        state <= 2'h0;
      end
    end
    hanning_signal_value <= _GEN_35[31:0];
  end
endmodule
module MyFifo(
  input         clock,
  input         reset,
  input  [31:0] io_datain_value,
  output [31:0] io_dataout_value,
  input         io_wr,
  input         io_rd,
  output        io_full,
  output        io_empty,
  output        io_MorethanN,
  output [31:0] io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_value [0:1023]; // @[Myfifo.scala 25:16]
  wire [31:0] mem_value__T_5_data; // @[Myfifo.scala 25:16]
  wire [9:0] mem_value__T_5_addr; // @[Myfifo.scala 25:16]
  wire [31:0] mem_value__T_33_data; // @[Myfifo.scala 25:16]
  wire [9:0] mem_value__T_33_addr; // @[Myfifo.scala 25:16]
  wire [31:0] mem_value__T_11_data; // @[Myfifo.scala 25:16]
  wire [9:0] mem_value__T_11_addr; // @[Myfifo.scala 25:16]
  wire  mem_value__T_11_mask; // @[Myfifo.scala 25:16]
  wire  mem_value__T_11_en; // @[Myfifo.scala 25:16]
  wire [31:0] mem_value__T_21_data; // @[Myfifo.scala 25:16]
  wire [9:0] mem_value__T_21_addr; // @[Myfifo.scala 25:16]
  wire  mem_value__T_21_mask; // @[Myfifo.scala 25:16]
  wire  mem_value__T_21_en; // @[Myfifo.scala 25:16]
  reg [31:0] count; // @[Myfifo.scala 24:22]
  reg [31:0] wp; // @[Myfifo.scala 26:19]
  reg [31:0] rp; // @[Myfifo.scala 27:19]
  wire  _T_2 = io_wr & io_rd; // @[Myfifo.scala 38:25]
  wire  _T_3 = count == 32'h0; // @[Myfifo.scala 39:16]
  wire  _T_7 = rp == 32'h3ff; // @[Myfifo.scala 33:16]
  wire [31:0] _T_9 = rp + 32'h1; // @[Myfifo.scala 34:34]
  wire  _T_13 = wp == 32'h3ff; // @[Myfifo.scala 33:16]
  wire [31:0] _T_15 = wp + 32'h1; // @[Myfifo.scala 34:34]
  wire [31:0] _GEN_2 = _T_3 ? $signed(io_datain_value) : $signed(mem_value__T_5_data); // @[Myfifo.scala 39:25]
  wire  _GEN_5 = _T_3 ? 1'h0 : 1'h1; // @[Myfifo.scala 39:25]
  wire  _T_17 = ~io_rd; // @[Myfifo.scala 46:42]
  wire  _T_18 = io_wr & _T_17; // @[Myfifo.scala 46:33]
  wire  _T_19 = count < 32'h400; // @[Myfifo.scala 48:16]
  wire [31:0] _T_27 = count + 32'h1; // @[Myfifo.scala 51:22]
  wire  _T_28 = ~io_wr; // @[Myfifo.scala 53:22]
  wire  _T_30 = _T_28 & io_rd; // @[Myfifo.scala 53:34]
  wire  _T_31 = count > 32'h0; // @[Myfifo.scala 54:16]
  wire [31:0] _T_39 = count - 32'h1; // @[Myfifo.scala 57:22]
  wire [31:0] _GEN_23 = _T_31 ? $signed(mem_value__T_33_data) : $signed(32'sh0); // @[Myfifo.scala 54:23]
  wire  _GEN_28 = _T_30 & _T_31; // @[Myfifo.scala 53:55]
  wire [31:0] _GEN_29 = _T_30 ? $signed(_GEN_23) : $signed(32'sh0); // @[Myfifo.scala 53:55]
  wire [31:0] _GEN_32 = _T_18 ? $signed(32'sh0) : $signed(_GEN_29); // @[Myfifo.scala 46:55]
  wire  _GEN_35 = _T_18 & _T_19; // @[Myfifo.scala 46:55]
  wire  _GEN_42 = _T_18 ? 1'h0 : _GEN_28; // @[Myfifo.scala 46:55]
  assign mem_value__T_5_addr = rp[9:0];
  assign mem_value__T_5_data = mem_value[mem_value__T_5_addr]; // @[Myfifo.scala 25:16]
  assign mem_value__T_33_addr = rp[9:0];
  assign mem_value__T_33_data = mem_value[mem_value__T_33_addr]; // @[Myfifo.scala 25:16]
  assign mem_value__T_11_data = io_datain_value;
  assign mem_value__T_11_addr = wp[9:0];
  assign mem_value__T_11_mask = 1'h1;
  assign mem_value__T_11_en = _T_2 & _GEN_5;
  assign mem_value__T_21_data = io_datain_value;
  assign mem_value__T_21_addr = wp[9:0];
  assign mem_value__T_21_mask = 1'h1;
  assign mem_value__T_21_en = _T_2 ? 1'h0 : _GEN_35;
  assign io_dataout_value = _T_2 ? $signed(_GEN_2) : $signed(_GEN_32); // @[Myfifo.scala 39:38 Myfifo.scala 41:20 Myfifo.scala 47:22 Myfifo.scala 55:18 Myfifo.scala 59:24 Myfifo.scala 62:22]
  assign io_full = 32'h400 == count; // @[Myfifo.scala 65:11]
  assign io_empty = count == 32'h0; // @[Myfifo.scala 66:12]
  assign io_MorethanN = count > 32'h200; // @[Myfifo.scala 67:16]
  assign io_count = count; // @[Myfifo.scala 68:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem_value[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wp = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rp = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem_value__T_11_en & mem_value__T_11_mask) begin
      mem_value[mem_value__T_11_addr] <= mem_value__T_11_data; // @[Myfifo.scala 25:16]
    end
    if(mem_value__T_21_en & mem_value__T_21_mask) begin
      mem_value[mem_value__T_21_addr] <= mem_value__T_21_data; // @[Myfifo.scala 25:16]
    end
    if (reset) begin
      count <= 32'h0;
    end else if (!(_T_2)) begin
      if (_T_18) begin
        if (_T_19) begin
          count <= _T_27;
        end
      end else if (_T_30) begin
        if (_T_31) begin
          count <= _T_39;
        end
      end
    end
    if (reset) begin
      wp <= 32'h0;
    end else if (_T_2) begin
      if (!(_T_3)) begin
        if (_T_13) begin
          wp <= 32'h0;
        end else begin
          wp <= _T_15;
        end
      end
    end else if (_T_18) begin
      if (_T_19) begin
        if (_T_13) begin
          wp <= 32'h0;
        end else begin
          wp <= _T_15;
        end
      end
    end
    if (reset) begin
      rp <= 32'h0;
    end else if (_T_2) begin
      if (!(_T_3)) begin
        if (_T_7) begin
          rp <= 32'h0;
        end else begin
          rp <= _T_9;
        end
      end
    end else if (!(_T_18)) begin
      if (_T_30) begin
        if (_T_31) begin
          if (_T_7) begin
            rp <= 32'h0;
          end else begin
            rp <= _T_9;
          end
        end
      end
    end
  end
endmodule
module HanningWithFIFO(
  input         clock,
  input         reset,
  output        io_signal_ready,
  input         io_signal_valid,
  input  [31:0] io_signal_bits_value,
  output        io_cosines_ready,
  input         io_cosines_valid,
  input  [31:0] io_cosines_bits_value,
  input         io_HanningSignal_ready,
  output        io_HanningSignal_valid,
  output [31:0] io_HanningSignal_bits_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  Hanningblock_clock; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_reset; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_io_signal_ready; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_io_signal_valid; // @[HanningWithFIFO.scala 19:37]
  wire [31:0] Hanningblock_io_signal_bits_value; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_io_cosines_ready; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_io_cosines_valid; // @[HanningWithFIFO.scala 19:37]
  wire [31:0] Hanningblock_io_cosines_bits_value; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_io_HanningSignal_ready; // @[HanningWithFIFO.scala 19:37]
  wire  Hanningblock_io_HanningSignal_valid; // @[HanningWithFIFO.scala 19:37]
  wire [31:0] Hanningblock_io_HanningSignal_bits_value; // @[HanningWithFIFO.scala 19:37]
  wire  HanningFIFO_clock; // @[HanningWithFIFO.scala 20:35]
  wire  HanningFIFO_reset; // @[HanningWithFIFO.scala 20:35]
  wire [31:0] HanningFIFO_io_datain_value; // @[HanningWithFIFO.scala 20:35]
  wire [31:0] HanningFIFO_io_dataout_value; // @[HanningWithFIFO.scala 20:35]
  wire  HanningFIFO_io_wr; // @[HanningWithFIFO.scala 20:35]
  wire  HanningFIFO_io_rd; // @[HanningWithFIFO.scala 20:35]
  wire  HanningFIFO_io_full; // @[HanningWithFIFO.scala 20:35]
  wire  HanningFIFO_io_empty; // @[HanningWithFIFO.scala 20:35]
  wire  HanningFIFO_io_MorethanN; // @[HanningWithFIFO.scala 20:35]
  wire [31:0] HanningFIFO_io_count; // @[HanningWithFIFO.scala 20:35]
  reg  BurstValid; // @[HanningWithFIFO.scala 22:27]
  reg [31:0] BurstReadCnt; // @[HanningWithFIFO.scala 23:29]
  wire  _T = BurstReadCnt < 32'h200; // @[HanningWithFIFO.scala 25:33]
  wire  _T_1 = BurstReadCnt > 32'h0; // @[HanningWithFIFO.scala 25:64]
  wire  BurstTransEn = _T & _T_1; // @[HanningWithFIFO.scala 25:48]
  wire  _T_3 = io_HanningSignal_ready & BurstValid; // @[HanningWithFIFO.scala 27:31]
  wire [31:0] _T_5 = BurstReadCnt + 32'h1; // @[HanningWithFIFO.scala 28:34]
  wire  _GEN_0 = HanningFIFO_io_MorethanN | BurstValid; // @[HanningWithFIFO.scala 35:36]
  Hanning Hanningblock ( // @[HanningWithFIFO.scala 19:37]
    .clock(Hanningblock_clock),
    .reset(Hanningblock_reset),
    .io_signal_ready(Hanningblock_io_signal_ready),
    .io_signal_valid(Hanningblock_io_signal_valid),
    .io_signal_bits_value(Hanningblock_io_signal_bits_value),
    .io_cosines_ready(Hanningblock_io_cosines_ready),
    .io_cosines_valid(Hanningblock_io_cosines_valid),
    .io_cosines_bits_value(Hanningblock_io_cosines_bits_value),
    .io_HanningSignal_ready(Hanningblock_io_HanningSignal_ready),
    .io_HanningSignal_valid(Hanningblock_io_HanningSignal_valid),
    .io_HanningSignal_bits_value(Hanningblock_io_HanningSignal_bits_value)
  );
  MyFifo HanningFIFO ( // @[HanningWithFIFO.scala 20:35]
    .clock(HanningFIFO_clock),
    .reset(HanningFIFO_reset),
    .io_datain_value(HanningFIFO_io_datain_value),
    .io_dataout_value(HanningFIFO_io_dataout_value),
    .io_wr(HanningFIFO_io_wr),
    .io_rd(HanningFIFO_io_rd),
    .io_full(HanningFIFO_io_full),
    .io_empty(HanningFIFO_io_empty),
    .io_MorethanN(HanningFIFO_io_MorethanN),
    .io_count(HanningFIFO_io_count)
  );
  assign io_signal_ready = Hanningblock_io_signal_ready; // @[HanningWithFIFO.scala 38:26]
  assign io_cosines_ready = Hanningblock_io_cosines_ready; // @[HanningWithFIFO.scala 39:27]
  assign io_HanningSignal_valid = BurstValid; // @[HanningWithFIFO.scala 41:26]
  assign io_HanningSignal_bits_value = HanningFIFO_io_dataout_value; // @[HanningWithFIFO.scala 42:26]
  assign Hanningblock_clock = clock;
  assign Hanningblock_reset = reset;
  assign Hanningblock_io_signal_valid = io_signal_valid; // @[HanningWithFIFO.scala 38:26]
  assign Hanningblock_io_signal_bits_value = io_signal_bits_value; // @[HanningWithFIFO.scala 38:26]
  assign Hanningblock_io_cosines_valid = io_cosines_valid; // @[HanningWithFIFO.scala 39:27]
  assign Hanningblock_io_cosines_bits_value = io_cosines_bits_value; // @[HanningWithFIFO.scala 39:27]
  assign Hanningblock_io_HanningSignal_ready = ~HanningFIFO_io_full; // @[HanningWithFIFO.scala 47:39]
  assign HanningFIFO_clock = clock;
  assign HanningFIFO_reset = reset;
  assign HanningFIFO_io_datain_value = Hanningblock_io_HanningSignal_bits_value; // @[HanningWithFIFO.scala 45:25]
  assign HanningFIFO_io_wr = Hanningblock_io_HanningSignal_valid; // @[HanningWithFIFO.scala 46:21]
  assign HanningFIFO_io_rd = BurstReadCnt != 32'h0; // @[HanningWithFIFO.scala 49:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  BurstValid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  BurstReadCnt = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      BurstValid <= 1'h0;
    end else if (_T_3) begin
      BurstValid <= 1'h0;
    end else if (!(BurstTransEn)) begin
      BurstValid <= _GEN_0;
    end
    if (reset) begin
      BurstReadCnt <= 32'h0;
    end else if (_T_3) begin
      BurstReadCnt <= _T_5;
    end else if (BurstTransEn) begin
      BurstReadCnt <= _T_5;
    end else begin
      BurstReadCnt <= 32'h0;
    end
  end
endmodule
module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 32:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 33:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 46:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 47:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 84:28]
  wire [63:0] _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 84:52]
  wire [63:0] _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 84:40]
  wire [63:0] _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 85:28]
  wire [63:0] _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 85:52]
  wire [63:0] _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 85:40]
  wire [47:0] _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 84:15]
  wire [47:0] _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 85:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 84:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 85:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 90:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 90:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 90:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 90:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 90:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 90:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 37:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 51:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 90:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 111:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 111:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 112:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 112:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 38:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 38:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 39:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 39:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 52:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 52:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 53:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 53:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 91:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 91:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 92:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 92:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 132:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 132:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 133:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 133:11]
endmodule
module FFT(
  input         clock,
  input         reset,
  input  [31:0] io_dIn_re,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid,
  output        io_busy
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 116:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 116:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 137:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 137:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 137:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 37:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 51:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 51:22]
  reg [9:0] cnt; // @[FFT.scala 63:20]
  wire  busy = cnt != 10'h0; // @[FFT.scala 64:18]
  wire  _T = io_din_valid | busy; // @[FFT.scala 65:21]
  wire  _T_1 = cnt == 10'h2ff; // @[FFT.scala 66:20]
  wire [9:0] _T_3 = cnt + 10'h1; // @[FFT.scala 66:67]
  wire [31:0] _GEN_2 = 8'h1 == cnt[7:0] ? $signed(32'shfffb) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3 = 8'h2 == cnt[7:0] ? $signed(32'shffec) : $signed(_GEN_2); // @[FFT.scala 52:18]
  wire [31:0] _GEN_4 = 8'h3 == cnt[7:0] ? $signed(32'shffd4) : $signed(_GEN_3); // @[FFT.scala 52:18]
  wire [31:0] _GEN_5 = 8'h4 == cnt[7:0] ? $signed(32'shffb1) : $signed(_GEN_4); // @[FFT.scala 52:18]
  wire [31:0] _GEN_6 = 8'h5 == cnt[7:0] ? $signed(32'shff85) : $signed(_GEN_5); // @[FFT.scala 52:18]
  wire [31:0] _GEN_7 = 8'h6 == cnt[7:0] ? $signed(32'shff4e) : $signed(_GEN_6); // @[FFT.scala 52:18]
  wire [31:0] _GEN_8 = 8'h7 == cnt[7:0] ? $signed(32'shff0e) : $signed(_GEN_7); // @[FFT.scala 52:18]
  wire [31:0] _GEN_9 = 8'h8 == cnt[7:0] ? $signed(32'shfec4) : $signed(_GEN_8); // @[FFT.scala 52:18]
  wire [31:0] _GEN_10 = 8'h9 == cnt[7:0] ? $signed(32'shfe71) : $signed(_GEN_9); // @[FFT.scala 52:18]
  wire [31:0] _GEN_11 = 8'ha == cnt[7:0] ? $signed(32'shfe13) : $signed(_GEN_10); // @[FFT.scala 52:18]
  wire [31:0] _GEN_12 = 8'hb == cnt[7:0] ? $signed(32'shfdac) : $signed(_GEN_11); // @[FFT.scala 52:18]
  wire [31:0] _GEN_13 = 8'hc == cnt[7:0] ? $signed(32'shfd3b) : $signed(_GEN_12); // @[FFT.scala 52:18]
  wire [31:0] _GEN_14 = 8'hd == cnt[7:0] ? $signed(32'shfcc0) : $signed(_GEN_13); // @[FFT.scala 52:18]
  wire [31:0] _GEN_15 = 8'he == cnt[7:0] ? $signed(32'shfc3b) : $signed(_GEN_14); // @[FFT.scala 52:18]
  wire [31:0] _GEN_16 = 8'hf == cnt[7:0] ? $signed(32'shfbad) : $signed(_GEN_15); // @[FFT.scala 52:18]
  wire [31:0] _GEN_17 = 8'h10 == cnt[7:0] ? $signed(32'shfb15) : $signed(_GEN_16); // @[FFT.scala 52:18]
  wire [31:0] _GEN_18 = 8'h11 == cnt[7:0] ? $signed(32'shfa73) : $signed(_GEN_17); // @[FFT.scala 52:18]
  wire [31:0] _GEN_19 = 8'h12 == cnt[7:0] ? $signed(32'shf9c8) : $signed(_GEN_18); // @[FFT.scala 52:18]
  wire [31:0] _GEN_20 = 8'h13 == cnt[7:0] ? $signed(32'shf913) : $signed(_GEN_19); // @[FFT.scala 52:18]
  wire [31:0] _GEN_21 = 8'h14 == cnt[7:0] ? $signed(32'shf854) : $signed(_GEN_20); // @[FFT.scala 52:18]
  wire [31:0] _GEN_22 = 8'h15 == cnt[7:0] ? $signed(32'shf78c) : $signed(_GEN_21); // @[FFT.scala 52:18]
  wire [31:0] _GEN_23 = 8'h16 == cnt[7:0] ? $signed(32'shf6ba) : $signed(_GEN_22); // @[FFT.scala 52:18]
  wire [31:0] _GEN_24 = 8'h17 == cnt[7:0] ? $signed(32'shf5df) : $signed(_GEN_23); // @[FFT.scala 52:18]
  wire [31:0] _GEN_25 = 8'h18 == cnt[7:0] ? $signed(32'shf4fa) : $signed(_GEN_24); // @[FFT.scala 52:18]
  wire [31:0] _GEN_26 = 8'h19 == cnt[7:0] ? $signed(32'shf40c) : $signed(_GEN_25); // @[FFT.scala 52:18]
  wire [31:0] _GEN_27 = 8'h1a == cnt[7:0] ? $signed(32'shf314) : $signed(_GEN_26); // @[FFT.scala 52:18]
  wire [31:0] _GEN_28 = 8'h1b == cnt[7:0] ? $signed(32'shf213) : $signed(_GEN_27); // @[FFT.scala 52:18]
  wire [31:0] _GEN_29 = 8'h1c == cnt[7:0] ? $signed(32'shf109) : $signed(_GEN_28); // @[FFT.scala 52:18]
  wire [31:0] _GEN_30 = 8'h1d == cnt[7:0] ? $signed(32'sheff5) : $signed(_GEN_29); // @[FFT.scala 52:18]
  wire [31:0] _GEN_31 = 8'h1e == cnt[7:0] ? $signed(32'sheed9) : $signed(_GEN_30); // @[FFT.scala 52:18]
  wire [31:0] _GEN_32 = 8'h1f == cnt[7:0] ? $signed(32'shedb3) : $signed(_GEN_31); // @[FFT.scala 52:18]
  wire [31:0] _GEN_33 = 8'h20 == cnt[7:0] ? $signed(32'shec83) : $signed(_GEN_32); // @[FFT.scala 52:18]
  wire [31:0] _GEN_34 = 8'h21 == cnt[7:0] ? $signed(32'sheb4b) : $signed(_GEN_33); // @[FFT.scala 52:18]
  wire [31:0] _GEN_35 = 8'h22 == cnt[7:0] ? $signed(32'shea0a) : $signed(_GEN_34); // @[FFT.scala 52:18]
  wire [31:0] _GEN_36 = 8'h23 == cnt[7:0] ? $signed(32'she8bf) : $signed(_GEN_35); // @[FFT.scala 52:18]
  wire [31:0] _GEN_37 = 8'h24 == cnt[7:0] ? $signed(32'she76c) : $signed(_GEN_36); // @[FFT.scala 52:18]
  wire [31:0] _GEN_38 = 8'h25 == cnt[7:0] ? $signed(32'she610) : $signed(_GEN_37); // @[FFT.scala 52:18]
  wire [31:0] _GEN_39 = 8'h26 == cnt[7:0] ? $signed(32'she4aa) : $signed(_GEN_38); // @[FFT.scala 52:18]
  wire [31:0] _GEN_40 = 8'h27 == cnt[7:0] ? $signed(32'she33c) : $signed(_GEN_39); // @[FFT.scala 52:18]
  wire [31:0] _GEN_41 = 8'h28 == cnt[7:0] ? $signed(32'she1c6) : $signed(_GEN_40); // @[FFT.scala 52:18]
  wire [31:0] _GEN_42 = 8'h29 == cnt[7:0] ? $signed(32'she046) : $signed(_GEN_41); // @[FFT.scala 52:18]
  wire [31:0] _GEN_43 = 8'h2a == cnt[7:0] ? $signed(32'shdebe) : $signed(_GEN_42); // @[FFT.scala 52:18]
  wire [31:0] _GEN_44 = 8'h2b == cnt[7:0] ? $signed(32'shdd2d) : $signed(_GEN_43); // @[FFT.scala 52:18]
  wire [31:0] _GEN_45 = 8'h2c == cnt[7:0] ? $signed(32'shdb94) : $signed(_GEN_44); // @[FFT.scala 52:18]
  wire [31:0] _GEN_46 = 8'h2d == cnt[7:0] ? $signed(32'shd9f2) : $signed(_GEN_45); // @[FFT.scala 52:18]
  wire [31:0] _GEN_47 = 8'h2e == cnt[7:0] ? $signed(32'shd848) : $signed(_GEN_46); // @[FFT.scala 52:18]
  wire [31:0] _GEN_48 = 8'h2f == cnt[7:0] ? $signed(32'shd696) : $signed(_GEN_47); // @[FFT.scala 52:18]
  wire [31:0] _GEN_49 = 8'h30 == cnt[7:0] ? $signed(32'shd4db) : $signed(_GEN_48); // @[FFT.scala 52:18]
  wire [31:0] _GEN_50 = 8'h31 == cnt[7:0] ? $signed(32'shd318) : $signed(_GEN_49); // @[FFT.scala 52:18]
  wire [31:0] _GEN_51 = 8'h32 == cnt[7:0] ? $signed(32'shd14d) : $signed(_GEN_50); // @[FFT.scala 52:18]
  wire [31:0] _GEN_52 = 8'h33 == cnt[7:0] ? $signed(32'shcf7a) : $signed(_GEN_51); // @[FFT.scala 52:18]
  wire [31:0] _GEN_53 = 8'h34 == cnt[7:0] ? $signed(32'shcd9f) : $signed(_GEN_52); // @[FFT.scala 52:18]
  wire [31:0] _GEN_54 = 8'h35 == cnt[7:0] ? $signed(32'shcbbc) : $signed(_GEN_53); // @[FFT.scala 52:18]
  wire [31:0] _GEN_55 = 8'h36 == cnt[7:0] ? $signed(32'shc9d1) : $signed(_GEN_54); // @[FFT.scala 52:18]
  wire [31:0] _GEN_56 = 8'h37 == cnt[7:0] ? $signed(32'shc7de) : $signed(_GEN_55); // @[FFT.scala 52:18]
  wire [31:0] _GEN_57 = 8'h38 == cnt[7:0] ? $signed(32'shc5e4) : $signed(_GEN_56); // @[FFT.scala 52:18]
  wire [31:0] _GEN_58 = 8'h39 == cnt[7:0] ? $signed(32'shc3e2) : $signed(_GEN_57); // @[FFT.scala 52:18]
  wire [31:0] _GEN_59 = 8'h3a == cnt[7:0] ? $signed(32'shc1d8) : $signed(_GEN_58); // @[FFT.scala 52:18]
  wire [31:0] _GEN_60 = 8'h3b == cnt[7:0] ? $signed(32'shbfc7) : $signed(_GEN_59); // @[FFT.scala 52:18]
  wire [31:0] _GEN_61 = 8'h3c == cnt[7:0] ? $signed(32'shbdaf) : $signed(_GEN_60); // @[FFT.scala 52:18]
  wire [31:0] _GEN_62 = 8'h3d == cnt[7:0] ? $signed(32'shbb8f) : $signed(_GEN_61); // @[FFT.scala 52:18]
  wire [31:0] _GEN_63 = 8'h3e == cnt[7:0] ? $signed(32'shb968) : $signed(_GEN_62); // @[FFT.scala 52:18]
  wire [31:0] _GEN_64 = 8'h3f == cnt[7:0] ? $signed(32'shb73a) : $signed(_GEN_63); // @[FFT.scala 52:18]
  wire [31:0] _GEN_65 = 8'h40 == cnt[7:0] ? $signed(32'shb505) : $signed(_GEN_64); // @[FFT.scala 52:18]
  wire [31:0] _GEN_66 = 8'h41 == cnt[7:0] ? $signed(32'shb2c9) : $signed(_GEN_65); // @[FFT.scala 52:18]
  wire [31:0] _GEN_67 = 8'h42 == cnt[7:0] ? $signed(32'shb086) : $signed(_GEN_66); // @[FFT.scala 52:18]
  wire [31:0] _GEN_68 = 8'h43 == cnt[7:0] ? $signed(32'shae3c) : $signed(_GEN_67); // @[FFT.scala 52:18]
  wire [31:0] _GEN_69 = 8'h44 == cnt[7:0] ? $signed(32'shabeb) : $signed(_GEN_68); // @[FFT.scala 52:18]
  wire [31:0] _GEN_70 = 8'h45 == cnt[7:0] ? $signed(32'sha994) : $signed(_GEN_69); // @[FFT.scala 52:18]
  wire [31:0] _GEN_71 = 8'h46 == cnt[7:0] ? $signed(32'sha736) : $signed(_GEN_70); // @[FFT.scala 52:18]
  wire [31:0] _GEN_72 = 8'h47 == cnt[7:0] ? $signed(32'sha4d2) : $signed(_GEN_71); // @[FFT.scala 52:18]
  wire [31:0] _GEN_73 = 8'h48 == cnt[7:0] ? $signed(32'sha268) : $signed(_GEN_72); // @[FFT.scala 52:18]
  wire [31:0] _GEN_74 = 8'h49 == cnt[7:0] ? $signed(32'sh9ff7) : $signed(_GEN_73); // @[FFT.scala 52:18]
  wire [31:0] _GEN_75 = 8'h4a == cnt[7:0] ? $signed(32'sh9d80) : $signed(_GEN_74); // @[FFT.scala 52:18]
  wire [31:0] _GEN_76 = 8'h4b == cnt[7:0] ? $signed(32'sh9b03) : $signed(_GEN_75); // @[FFT.scala 52:18]
  wire [31:0] _GEN_77 = 8'h4c == cnt[7:0] ? $signed(32'sh9880) : $signed(_GEN_76); // @[FFT.scala 52:18]
  wire [31:0] _GEN_78 = 8'h4d == cnt[7:0] ? $signed(32'sh95f7) : $signed(_GEN_77); // @[FFT.scala 52:18]
  wire [31:0] _GEN_79 = 8'h4e == cnt[7:0] ? $signed(32'sh9368) : $signed(_GEN_78); // @[FFT.scala 52:18]
  wire [31:0] _GEN_80 = 8'h4f == cnt[7:0] ? $signed(32'sh90d4) : $signed(_GEN_79); // @[FFT.scala 52:18]
  wire [31:0] _GEN_81 = 8'h50 == cnt[7:0] ? $signed(32'sh8e3a) : $signed(_GEN_80); // @[FFT.scala 52:18]
  wire [31:0] _GEN_82 = 8'h51 == cnt[7:0] ? $signed(32'sh8b9a) : $signed(_GEN_81); // @[FFT.scala 52:18]
  wire [31:0] _GEN_83 = 8'h52 == cnt[7:0] ? $signed(32'sh88f6) : $signed(_GEN_82); // @[FFT.scala 52:18]
  wire [31:0] _GEN_84 = 8'h53 == cnt[7:0] ? $signed(32'sh864c) : $signed(_GEN_83); // @[FFT.scala 52:18]
  wire [31:0] _GEN_85 = 8'h54 == cnt[7:0] ? $signed(32'sh839c) : $signed(_GEN_84); // @[FFT.scala 52:18]
  wire [31:0] _GEN_86 = 8'h55 == cnt[7:0] ? $signed(32'sh80e8) : $signed(_GEN_85); // @[FFT.scala 52:18]
  wire [31:0] _GEN_87 = 8'h56 == cnt[7:0] ? $signed(32'sh7e2f) : $signed(_GEN_86); // @[FFT.scala 52:18]
  wire [31:0] _GEN_88 = 8'h57 == cnt[7:0] ? $signed(32'sh7b70) : $signed(_GEN_87); // @[FFT.scala 52:18]
  wire [31:0] _GEN_89 = 8'h58 == cnt[7:0] ? $signed(32'sh78ad) : $signed(_GEN_88); // @[FFT.scala 52:18]
  wire [31:0] _GEN_90 = 8'h59 == cnt[7:0] ? $signed(32'sh75e6) : $signed(_GEN_89); // @[FFT.scala 52:18]
  wire [31:0] _GEN_91 = 8'h5a == cnt[7:0] ? $signed(32'sh731a) : $signed(_GEN_90); // @[FFT.scala 52:18]
  wire [31:0] _GEN_92 = 8'h5b == cnt[7:0] ? $signed(32'sh7049) : $signed(_GEN_91); // @[FFT.scala 52:18]
  wire [31:0] _GEN_93 = 8'h5c == cnt[7:0] ? $signed(32'sh6d74) : $signed(_GEN_92); // @[FFT.scala 52:18]
  wire [31:0] _GEN_94 = 8'h5d == cnt[7:0] ? $signed(32'sh6a9b) : $signed(_GEN_93); // @[FFT.scala 52:18]
  wire [31:0] _GEN_95 = 8'h5e == cnt[7:0] ? $signed(32'sh67be) : $signed(_GEN_94); // @[FFT.scala 52:18]
  wire [31:0] _GEN_96 = 8'h5f == cnt[7:0] ? $signed(32'sh64dd) : $signed(_GEN_95); // @[FFT.scala 52:18]
  wire [31:0] _GEN_97 = 8'h60 == cnt[7:0] ? $signed(32'sh61f8) : $signed(_GEN_96); // @[FFT.scala 52:18]
  wire [31:0] _GEN_98 = 8'h61 == cnt[7:0] ? $signed(32'sh5f0f) : $signed(_GEN_97); // @[FFT.scala 52:18]
  wire [31:0] _GEN_99 = 8'h62 == cnt[7:0] ? $signed(32'sh5c22) : $signed(_GEN_98); // @[FFT.scala 52:18]
  wire [31:0] _GEN_100 = 8'h63 == cnt[7:0] ? $signed(32'sh5932) : $signed(_GEN_99); // @[FFT.scala 52:18]
  wire [31:0] _GEN_101 = 8'h64 == cnt[7:0] ? $signed(32'sh563e) : $signed(_GEN_100); // @[FFT.scala 52:18]
  wire [31:0] _GEN_102 = 8'h65 == cnt[7:0] ? $signed(32'sh5348) : $signed(_GEN_101); // @[FFT.scala 52:18]
  wire [31:0] _GEN_103 = 8'h66 == cnt[7:0] ? $signed(32'sh504d) : $signed(_GEN_102); // @[FFT.scala 52:18]
  wire [31:0] _GEN_104 = 8'h67 == cnt[7:0] ? $signed(32'sh4d50) : $signed(_GEN_103); // @[FFT.scala 52:18]
  wire [31:0] _GEN_105 = 8'h68 == cnt[7:0] ? $signed(32'sh4a50) : $signed(_GEN_104); // @[FFT.scala 52:18]
  wire [31:0] _GEN_106 = 8'h69 == cnt[7:0] ? $signed(32'sh474d) : $signed(_GEN_105); // @[FFT.scala 52:18]
  wire [31:0] _GEN_107 = 8'h6a == cnt[7:0] ? $signed(32'sh4447) : $signed(_GEN_106); // @[FFT.scala 52:18]
  wire [31:0] _GEN_108 = 8'h6b == cnt[7:0] ? $signed(32'sh413f) : $signed(_GEN_107); // @[FFT.scala 52:18]
  wire [31:0] _GEN_109 = 8'h6c == cnt[7:0] ? $signed(32'sh3e34) : $signed(_GEN_108); // @[FFT.scala 52:18]
  wire [31:0] _GEN_110 = 8'h6d == cnt[7:0] ? $signed(32'sh3b27) : $signed(_GEN_109); // @[FFT.scala 52:18]
  wire [31:0] _GEN_111 = 8'h6e == cnt[7:0] ? $signed(32'sh3817) : $signed(_GEN_110); // @[FFT.scala 52:18]
  wire [31:0] _GEN_112 = 8'h6f == cnt[7:0] ? $signed(32'sh3505) : $signed(_GEN_111); // @[FFT.scala 52:18]
  wire [31:0] _GEN_113 = 8'h70 == cnt[7:0] ? $signed(32'sh31f1) : $signed(_GEN_112); // @[FFT.scala 52:18]
  wire [31:0] _GEN_114 = 8'h71 == cnt[7:0] ? $signed(32'sh2edc) : $signed(_GEN_113); // @[FFT.scala 52:18]
  wire [31:0] _GEN_115 = 8'h72 == cnt[7:0] ? $signed(32'sh2bc4) : $signed(_GEN_114); // @[FFT.scala 52:18]
  wire [31:0] _GEN_116 = 8'h73 == cnt[7:0] ? $signed(32'sh28ab) : $signed(_GEN_115); // @[FFT.scala 52:18]
  wire [31:0] _GEN_117 = 8'h74 == cnt[7:0] ? $signed(32'sh2590) : $signed(_GEN_116); // @[FFT.scala 52:18]
  wire [31:0] _GEN_118 = 8'h75 == cnt[7:0] ? $signed(32'sh2274) : $signed(_GEN_117); // @[FFT.scala 52:18]
  wire [31:0] _GEN_119 = 8'h76 == cnt[7:0] ? $signed(32'sh1f56) : $signed(_GEN_118); // @[FFT.scala 52:18]
  wire [31:0] _GEN_120 = 8'h77 == cnt[7:0] ? $signed(32'sh1c38) : $signed(_GEN_119); // @[FFT.scala 52:18]
  wire [31:0] _GEN_121 = 8'h78 == cnt[7:0] ? $signed(32'sh1918) : $signed(_GEN_120); // @[FFT.scala 52:18]
  wire [31:0] _GEN_122 = 8'h79 == cnt[7:0] ? $signed(32'sh15f7) : $signed(_GEN_121); // @[FFT.scala 52:18]
  wire [31:0] _GEN_123 = 8'h7a == cnt[7:0] ? $signed(32'sh12d5) : $signed(_GEN_122); // @[FFT.scala 52:18]
  wire [31:0] _GEN_124 = 8'h7b == cnt[7:0] ? $signed(32'shfb3) : $signed(_GEN_123); // @[FFT.scala 52:18]
  wire [31:0] _GEN_125 = 8'h7c == cnt[7:0] ? $signed(32'shc90) : $signed(_GEN_124); // @[FFT.scala 52:18]
  wire [31:0] _GEN_126 = 8'h7d == cnt[7:0] ? $signed(32'sh96c) : $signed(_GEN_125); // @[FFT.scala 52:18]
  wire [31:0] _GEN_127 = 8'h7e == cnt[7:0] ? $signed(32'sh648) : $signed(_GEN_126); // @[FFT.scala 52:18]
  wire [31:0] _GEN_128 = 8'h7f == cnt[7:0] ? $signed(32'sh324) : $signed(_GEN_127); // @[FFT.scala 52:18]
  wire [31:0] _GEN_129 = 8'h80 == cnt[7:0] ? $signed(32'sh0) : $signed(_GEN_128); // @[FFT.scala 52:18]
  wire [31:0] _GEN_130 = 8'h81 == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_129); // @[FFT.scala 52:18]
  wire [31:0] _GEN_131 = 8'h82 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_130); // @[FFT.scala 52:18]
  wire [31:0] _GEN_132 = 8'h83 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_131); // @[FFT.scala 52:18]
  wire [31:0] _GEN_133 = 8'h84 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_132); // @[FFT.scala 52:18]
  wire [31:0] _GEN_134 = 8'h85 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_133); // @[FFT.scala 52:18]
  wire [31:0] _GEN_135 = 8'h86 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_134); // @[FFT.scala 52:18]
  wire [31:0] _GEN_136 = 8'h87 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_135); // @[FFT.scala 52:18]
  wire [31:0] _GEN_137 = 8'h88 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_136); // @[FFT.scala 52:18]
  wire [31:0] _GEN_138 = 8'h89 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_137); // @[FFT.scala 52:18]
  wire [31:0] _GEN_139 = 8'h8a == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_138); // @[FFT.scala 52:18]
  wire [31:0] _GEN_140 = 8'h8b == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_139); // @[FFT.scala 52:18]
  wire [31:0] _GEN_141 = 8'h8c == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_140); // @[FFT.scala 52:18]
  wire [31:0] _GEN_142 = 8'h8d == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_141); // @[FFT.scala 52:18]
  wire [31:0] _GEN_143 = 8'h8e == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_142); // @[FFT.scala 52:18]
  wire [31:0] _GEN_144 = 8'h8f == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_143); // @[FFT.scala 52:18]
  wire [31:0] _GEN_145 = 8'h90 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_144); // @[FFT.scala 52:18]
  wire [31:0] _GEN_146 = 8'h91 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_145); // @[FFT.scala 52:18]
  wire [31:0] _GEN_147 = 8'h92 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_146); // @[FFT.scala 52:18]
  wire [31:0] _GEN_148 = 8'h93 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_147); // @[FFT.scala 52:18]
  wire [31:0] _GEN_149 = 8'h94 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_148); // @[FFT.scala 52:18]
  wire [31:0] _GEN_150 = 8'h95 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_149); // @[FFT.scala 52:18]
  wire [31:0] _GEN_151 = 8'h96 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_150); // @[FFT.scala 52:18]
  wire [31:0] _GEN_152 = 8'h97 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_151); // @[FFT.scala 52:18]
  wire [31:0] _GEN_153 = 8'h98 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_152); // @[FFT.scala 52:18]
  wire [31:0] _GEN_154 = 8'h99 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_153); // @[FFT.scala 52:18]
  wire [31:0] _GEN_155 = 8'h9a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_154); // @[FFT.scala 52:18]
  wire [31:0] _GEN_156 = 8'h9b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_155); // @[FFT.scala 52:18]
  wire [31:0] _GEN_157 = 8'h9c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_156); // @[FFT.scala 52:18]
  wire [31:0] _GEN_158 = 8'h9d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_157); // @[FFT.scala 52:18]
  wire [31:0] _GEN_159 = 8'h9e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_158); // @[FFT.scala 52:18]
  wire [31:0] _GEN_160 = 8'h9f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_159); // @[FFT.scala 52:18]
  wire [31:0] _GEN_161 = 8'ha0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_160); // @[FFT.scala 52:18]
  wire [31:0] _GEN_162 = 8'ha1 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_161); // @[FFT.scala 52:18]
  wire [31:0] _GEN_163 = 8'ha2 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_162); // @[FFT.scala 52:18]
  wire [31:0] _GEN_164 = 8'ha3 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_163); // @[FFT.scala 52:18]
  wire [31:0] _GEN_165 = 8'ha4 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_164); // @[FFT.scala 52:18]
  wire [31:0] _GEN_166 = 8'ha5 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_165); // @[FFT.scala 52:18]
  wire [31:0] _GEN_167 = 8'ha6 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_166); // @[FFT.scala 52:18]
  wire [31:0] _GEN_168 = 8'ha7 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_167); // @[FFT.scala 52:18]
  wire [31:0] _GEN_169 = 8'ha8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_168); // @[FFT.scala 52:18]
  wire [31:0] _GEN_170 = 8'ha9 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_169); // @[FFT.scala 52:18]
  wire [31:0] _GEN_171 = 8'haa == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_170); // @[FFT.scala 52:18]
  wire [31:0] _GEN_172 = 8'hab == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_171); // @[FFT.scala 52:18]
  wire [31:0] _GEN_173 = 8'hac == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_172); // @[FFT.scala 52:18]
  wire [31:0] _GEN_174 = 8'had == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_173); // @[FFT.scala 52:18]
  wire [31:0] _GEN_175 = 8'hae == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_174); // @[FFT.scala 52:18]
  wire [31:0] _GEN_176 = 8'haf == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_175); // @[FFT.scala 52:18]
  wire [31:0] _GEN_177 = 8'hb0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_176); // @[FFT.scala 52:18]
  wire [31:0] _GEN_178 = 8'hb1 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_177); // @[FFT.scala 52:18]
  wire [31:0] _GEN_179 = 8'hb2 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_178); // @[FFT.scala 52:18]
  wire [31:0] _GEN_180 = 8'hb3 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_179); // @[FFT.scala 52:18]
  wire [31:0] _GEN_181 = 8'hb4 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_180); // @[FFT.scala 52:18]
  wire [31:0] _GEN_182 = 8'hb5 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_181); // @[FFT.scala 52:18]
  wire [31:0] _GEN_183 = 8'hb6 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_182); // @[FFT.scala 52:18]
  wire [31:0] _GEN_184 = 8'hb7 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_183); // @[FFT.scala 52:18]
  wire [31:0] _GEN_185 = 8'hb8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_184); // @[FFT.scala 52:18]
  wire [31:0] _GEN_186 = 8'hb9 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_185); // @[FFT.scala 52:18]
  wire [31:0] _GEN_187 = 8'hba == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_186); // @[FFT.scala 52:18]
  wire [31:0] _GEN_188 = 8'hbb == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_187); // @[FFT.scala 52:18]
  wire [31:0] _GEN_189 = 8'hbc == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_188); // @[FFT.scala 52:18]
  wire [31:0] _GEN_190 = 8'hbd == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_189); // @[FFT.scala 52:18]
  wire [31:0] _GEN_191 = 8'hbe == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_190); // @[FFT.scala 52:18]
  wire [31:0] _GEN_192 = 8'hbf == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_191); // @[FFT.scala 52:18]
  wire [31:0] _GEN_193 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_192); // @[FFT.scala 52:18]
  wire [31:0] _GEN_194 = 8'hc1 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_193); // @[FFT.scala 52:18]
  wire [31:0] _GEN_195 = 8'hc2 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_194); // @[FFT.scala 52:18]
  wire [31:0] _GEN_196 = 8'hc3 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_195); // @[FFT.scala 52:18]
  wire [31:0] _GEN_197 = 8'hc4 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_196); // @[FFT.scala 52:18]
  wire [31:0] _GEN_198 = 8'hc5 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_197); // @[FFT.scala 52:18]
  wire [31:0] _GEN_199 = 8'hc6 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_198); // @[FFT.scala 52:18]
  wire [31:0] _GEN_200 = 8'hc7 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_199); // @[FFT.scala 52:18]
  wire [31:0] _GEN_201 = 8'hc8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_200); // @[FFT.scala 52:18]
  wire [31:0] _GEN_202 = 8'hc9 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_201); // @[FFT.scala 52:18]
  wire [31:0] _GEN_203 = 8'hca == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_202); // @[FFT.scala 52:18]
  wire [31:0] _GEN_204 = 8'hcb == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_203); // @[FFT.scala 52:18]
  wire [31:0] _GEN_205 = 8'hcc == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_204); // @[FFT.scala 52:18]
  wire [31:0] _GEN_206 = 8'hcd == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_205); // @[FFT.scala 52:18]
  wire [31:0] _GEN_207 = 8'hce == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_206); // @[FFT.scala 52:18]
  wire [31:0] _GEN_208 = 8'hcf == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_207); // @[FFT.scala 52:18]
  wire [31:0] _GEN_209 = 8'hd0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_208); // @[FFT.scala 52:18]
  wire [31:0] _GEN_210 = 8'hd1 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_209); // @[FFT.scala 52:18]
  wire [31:0] _GEN_211 = 8'hd2 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_210); // @[FFT.scala 52:18]
  wire [31:0] _GEN_212 = 8'hd3 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_211); // @[FFT.scala 52:18]
  wire [31:0] _GEN_213 = 8'hd4 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_212); // @[FFT.scala 52:18]
  wire [31:0] _GEN_214 = 8'hd5 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_213); // @[FFT.scala 52:18]
  wire [31:0] _GEN_215 = 8'hd6 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_214); // @[FFT.scala 52:18]
  wire [31:0] _GEN_216 = 8'hd7 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_215); // @[FFT.scala 52:18]
  wire [31:0] _GEN_217 = 8'hd8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_216); // @[FFT.scala 52:18]
  wire [31:0] _GEN_218 = 8'hd9 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_217); // @[FFT.scala 52:18]
  wire [31:0] _GEN_219 = 8'hda == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_218); // @[FFT.scala 52:18]
  wire [31:0] _GEN_220 = 8'hdb == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_219); // @[FFT.scala 52:18]
  wire [31:0] _GEN_221 = 8'hdc == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_220); // @[FFT.scala 52:18]
  wire [31:0] _GEN_222 = 8'hdd == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_221); // @[FFT.scala 52:18]
  wire [31:0] _GEN_223 = 8'hde == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_222); // @[FFT.scala 52:18]
  wire [31:0] _GEN_224 = 8'hdf == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_223); // @[FFT.scala 52:18]
  wire [31:0] _GEN_225 = 8'he0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_224); // @[FFT.scala 52:18]
  wire [31:0] _GEN_226 = 8'he1 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_225); // @[FFT.scala 52:18]
  wire [31:0] _GEN_227 = 8'he2 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_226); // @[FFT.scala 52:18]
  wire [31:0] _GEN_228 = 8'he3 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_227); // @[FFT.scala 52:18]
  wire [31:0] _GEN_229 = 8'he4 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_228); // @[FFT.scala 52:18]
  wire [31:0] _GEN_230 = 8'he5 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_229); // @[FFT.scala 52:18]
  wire [31:0] _GEN_231 = 8'he6 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_230); // @[FFT.scala 52:18]
  wire [31:0] _GEN_232 = 8'he7 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_231); // @[FFT.scala 52:18]
  wire [31:0] _GEN_233 = 8'he8 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_232); // @[FFT.scala 52:18]
  wire [31:0] _GEN_234 = 8'he9 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_233); // @[FFT.scala 52:18]
  wire [31:0] _GEN_235 = 8'hea == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_234); // @[FFT.scala 52:18]
  wire [31:0] _GEN_236 = 8'heb == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_235); // @[FFT.scala 52:18]
  wire [31:0] _GEN_237 = 8'hec == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_236); // @[FFT.scala 52:18]
  wire [31:0] _GEN_238 = 8'hed == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_237); // @[FFT.scala 52:18]
  wire [31:0] _GEN_239 = 8'hee == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_238); // @[FFT.scala 52:18]
  wire [31:0] _GEN_240 = 8'hef == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_239); // @[FFT.scala 52:18]
  wire [31:0] _GEN_241 = 8'hf0 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_240); // @[FFT.scala 52:18]
  wire [31:0] _GEN_242 = 8'hf1 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_241); // @[FFT.scala 52:18]
  wire [31:0] _GEN_243 = 8'hf2 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_242); // @[FFT.scala 52:18]
  wire [31:0] _GEN_244 = 8'hf3 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_243); // @[FFT.scala 52:18]
  wire [31:0] _GEN_245 = 8'hf4 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_244); // @[FFT.scala 52:18]
  wire [31:0] _GEN_246 = 8'hf5 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_245); // @[FFT.scala 52:18]
  wire [31:0] _GEN_247 = 8'hf6 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_246); // @[FFT.scala 52:18]
  wire [31:0] _GEN_248 = 8'hf7 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_247); // @[FFT.scala 52:18]
  wire [31:0] _GEN_249 = 8'hf8 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_248); // @[FFT.scala 52:18]
  wire [31:0] _GEN_250 = 8'hf9 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_249); // @[FFT.scala 52:18]
  wire [31:0] _GEN_251 = 8'hfa == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_250); // @[FFT.scala 52:18]
  wire [31:0] _GEN_252 = 8'hfb == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_251); // @[FFT.scala 52:18]
  wire [31:0] _GEN_253 = 8'hfc == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_252); // @[FFT.scala 52:18]
  wire [31:0] _GEN_254 = 8'hfd == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_253); // @[FFT.scala 52:18]
  wire [31:0] _GEN_255 = 8'hfe == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_254); // @[FFT.scala 52:18]
  wire [31:0] _GEN_770 = 8'h1 == cnt[7:0] ? $signed(-32'sh324) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_771 = 8'h2 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_770); // @[FFT.scala 53:18]
  wire [31:0] _GEN_772 = 8'h3 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_771); // @[FFT.scala 53:18]
  wire [31:0] _GEN_773 = 8'h4 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_772); // @[FFT.scala 53:18]
  wire [31:0] _GEN_774 = 8'h5 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_773); // @[FFT.scala 53:18]
  wire [31:0] _GEN_775 = 8'h6 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_774); // @[FFT.scala 53:18]
  wire [31:0] _GEN_776 = 8'h7 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_775); // @[FFT.scala 53:18]
  wire [31:0] _GEN_777 = 8'h8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_776); // @[FFT.scala 53:18]
  wire [31:0] _GEN_778 = 8'h9 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_777); // @[FFT.scala 53:18]
  wire [31:0] _GEN_779 = 8'ha == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_778); // @[FFT.scala 53:18]
  wire [31:0] _GEN_780 = 8'hb == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_779); // @[FFT.scala 53:18]
  wire [31:0] _GEN_781 = 8'hc == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_780); // @[FFT.scala 53:18]
  wire [31:0] _GEN_782 = 8'hd == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_781); // @[FFT.scala 53:18]
  wire [31:0] _GEN_783 = 8'he == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_782); // @[FFT.scala 53:18]
  wire [31:0] _GEN_784 = 8'hf == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_783); // @[FFT.scala 53:18]
  wire [31:0] _GEN_785 = 8'h10 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_784); // @[FFT.scala 53:18]
  wire [31:0] _GEN_786 = 8'h11 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_785); // @[FFT.scala 53:18]
  wire [31:0] _GEN_787 = 8'h12 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_786); // @[FFT.scala 53:18]
  wire [31:0] _GEN_788 = 8'h13 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_787); // @[FFT.scala 53:18]
  wire [31:0] _GEN_789 = 8'h14 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_788); // @[FFT.scala 53:18]
  wire [31:0] _GEN_790 = 8'h15 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_789); // @[FFT.scala 53:18]
  wire [31:0] _GEN_791 = 8'h16 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_790); // @[FFT.scala 53:18]
  wire [31:0] _GEN_792 = 8'h17 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_791); // @[FFT.scala 53:18]
  wire [31:0] _GEN_793 = 8'h18 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_792); // @[FFT.scala 53:18]
  wire [31:0] _GEN_794 = 8'h19 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_793); // @[FFT.scala 53:18]
  wire [31:0] _GEN_795 = 8'h1a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_794); // @[FFT.scala 53:18]
  wire [31:0] _GEN_796 = 8'h1b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_795); // @[FFT.scala 53:18]
  wire [31:0] _GEN_797 = 8'h1c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_796); // @[FFT.scala 53:18]
  wire [31:0] _GEN_798 = 8'h1d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_797); // @[FFT.scala 53:18]
  wire [31:0] _GEN_799 = 8'h1e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_798); // @[FFT.scala 53:18]
  wire [31:0] _GEN_800 = 8'h1f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_799); // @[FFT.scala 53:18]
  wire [31:0] _GEN_801 = 8'h20 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_800); // @[FFT.scala 53:18]
  wire [31:0] _GEN_802 = 8'h21 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_801); // @[FFT.scala 53:18]
  wire [31:0] _GEN_803 = 8'h22 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_802); // @[FFT.scala 53:18]
  wire [31:0] _GEN_804 = 8'h23 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_803); // @[FFT.scala 53:18]
  wire [31:0] _GEN_805 = 8'h24 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_804); // @[FFT.scala 53:18]
  wire [31:0] _GEN_806 = 8'h25 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_805); // @[FFT.scala 53:18]
  wire [31:0] _GEN_807 = 8'h26 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_806); // @[FFT.scala 53:18]
  wire [31:0] _GEN_808 = 8'h27 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_807); // @[FFT.scala 53:18]
  wire [31:0] _GEN_809 = 8'h28 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_808); // @[FFT.scala 53:18]
  wire [31:0] _GEN_810 = 8'h29 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_809); // @[FFT.scala 53:18]
  wire [31:0] _GEN_811 = 8'h2a == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_810); // @[FFT.scala 53:18]
  wire [31:0] _GEN_812 = 8'h2b == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_811); // @[FFT.scala 53:18]
  wire [31:0] _GEN_813 = 8'h2c == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_812); // @[FFT.scala 53:18]
  wire [31:0] _GEN_814 = 8'h2d == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_813); // @[FFT.scala 53:18]
  wire [31:0] _GEN_815 = 8'h2e == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_814); // @[FFT.scala 53:18]
  wire [31:0] _GEN_816 = 8'h2f == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_815); // @[FFT.scala 53:18]
  wire [31:0] _GEN_817 = 8'h30 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_816); // @[FFT.scala 53:18]
  wire [31:0] _GEN_818 = 8'h31 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_817); // @[FFT.scala 53:18]
  wire [31:0] _GEN_819 = 8'h32 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_818); // @[FFT.scala 53:18]
  wire [31:0] _GEN_820 = 8'h33 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_819); // @[FFT.scala 53:18]
  wire [31:0] _GEN_821 = 8'h34 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_820); // @[FFT.scala 53:18]
  wire [31:0] _GEN_822 = 8'h35 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_821); // @[FFT.scala 53:18]
  wire [31:0] _GEN_823 = 8'h36 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_822); // @[FFT.scala 53:18]
  wire [31:0] _GEN_824 = 8'h37 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_823); // @[FFT.scala 53:18]
  wire [31:0] _GEN_825 = 8'h38 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_824); // @[FFT.scala 53:18]
  wire [31:0] _GEN_826 = 8'h39 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_825); // @[FFT.scala 53:18]
  wire [31:0] _GEN_827 = 8'h3a == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_826); // @[FFT.scala 53:18]
  wire [31:0] _GEN_828 = 8'h3b == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_827); // @[FFT.scala 53:18]
  wire [31:0] _GEN_829 = 8'h3c == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_828); // @[FFT.scala 53:18]
  wire [31:0] _GEN_830 = 8'h3d == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_829); // @[FFT.scala 53:18]
  wire [31:0] _GEN_831 = 8'h3e == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_830); // @[FFT.scala 53:18]
  wire [31:0] _GEN_832 = 8'h3f == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_831); // @[FFT.scala 53:18]
  wire [31:0] _GEN_833 = 8'h40 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_832); // @[FFT.scala 53:18]
  wire [31:0] _GEN_834 = 8'h41 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_833); // @[FFT.scala 53:18]
  wire [31:0] _GEN_835 = 8'h42 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_834); // @[FFT.scala 53:18]
  wire [31:0] _GEN_836 = 8'h43 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_835); // @[FFT.scala 53:18]
  wire [31:0] _GEN_837 = 8'h44 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_836); // @[FFT.scala 53:18]
  wire [31:0] _GEN_838 = 8'h45 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_837); // @[FFT.scala 53:18]
  wire [31:0] _GEN_839 = 8'h46 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_838); // @[FFT.scala 53:18]
  wire [31:0] _GEN_840 = 8'h47 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_839); // @[FFT.scala 53:18]
  wire [31:0] _GEN_841 = 8'h48 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_840); // @[FFT.scala 53:18]
  wire [31:0] _GEN_842 = 8'h49 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_841); // @[FFT.scala 53:18]
  wire [31:0] _GEN_843 = 8'h4a == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_842); // @[FFT.scala 53:18]
  wire [31:0] _GEN_844 = 8'h4b == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_843); // @[FFT.scala 53:18]
  wire [31:0] _GEN_845 = 8'h4c == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_844); // @[FFT.scala 53:18]
  wire [31:0] _GEN_846 = 8'h4d == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_845); // @[FFT.scala 53:18]
  wire [31:0] _GEN_847 = 8'h4e == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_846); // @[FFT.scala 53:18]
  wire [31:0] _GEN_848 = 8'h4f == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_847); // @[FFT.scala 53:18]
  wire [31:0] _GEN_849 = 8'h50 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_848); // @[FFT.scala 53:18]
  wire [31:0] _GEN_850 = 8'h51 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_849); // @[FFT.scala 53:18]
  wire [31:0] _GEN_851 = 8'h52 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_850); // @[FFT.scala 53:18]
  wire [31:0] _GEN_852 = 8'h53 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_851); // @[FFT.scala 53:18]
  wire [31:0] _GEN_853 = 8'h54 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_852); // @[FFT.scala 53:18]
  wire [31:0] _GEN_854 = 8'h55 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_853); // @[FFT.scala 53:18]
  wire [31:0] _GEN_855 = 8'h56 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_854); // @[FFT.scala 53:18]
  wire [31:0] _GEN_856 = 8'h57 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_855); // @[FFT.scala 53:18]
  wire [31:0] _GEN_857 = 8'h58 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_856); // @[FFT.scala 53:18]
  wire [31:0] _GEN_858 = 8'h59 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_857); // @[FFT.scala 53:18]
  wire [31:0] _GEN_859 = 8'h5a == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_858); // @[FFT.scala 53:18]
  wire [31:0] _GEN_860 = 8'h5b == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_859); // @[FFT.scala 53:18]
  wire [31:0] _GEN_861 = 8'h5c == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_860); // @[FFT.scala 53:18]
  wire [31:0] _GEN_862 = 8'h5d == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_861); // @[FFT.scala 53:18]
  wire [31:0] _GEN_863 = 8'h5e == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_862); // @[FFT.scala 53:18]
  wire [31:0] _GEN_864 = 8'h5f == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_863); // @[FFT.scala 53:18]
  wire [31:0] _GEN_865 = 8'h60 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_864); // @[FFT.scala 53:18]
  wire [31:0] _GEN_866 = 8'h61 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_865); // @[FFT.scala 53:18]
  wire [31:0] _GEN_867 = 8'h62 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_866); // @[FFT.scala 53:18]
  wire [31:0] _GEN_868 = 8'h63 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_867); // @[FFT.scala 53:18]
  wire [31:0] _GEN_869 = 8'h64 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_868); // @[FFT.scala 53:18]
  wire [31:0] _GEN_870 = 8'h65 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_869); // @[FFT.scala 53:18]
  wire [31:0] _GEN_871 = 8'h66 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_870); // @[FFT.scala 53:18]
  wire [31:0] _GEN_872 = 8'h67 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_871); // @[FFT.scala 53:18]
  wire [31:0] _GEN_873 = 8'h68 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_872); // @[FFT.scala 53:18]
  wire [31:0] _GEN_874 = 8'h69 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_873); // @[FFT.scala 53:18]
  wire [31:0] _GEN_875 = 8'h6a == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_874); // @[FFT.scala 53:18]
  wire [31:0] _GEN_876 = 8'h6b == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_875); // @[FFT.scala 53:18]
  wire [31:0] _GEN_877 = 8'h6c == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_876); // @[FFT.scala 53:18]
  wire [31:0] _GEN_878 = 8'h6d == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_877); // @[FFT.scala 53:18]
  wire [31:0] _GEN_879 = 8'h6e == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_878); // @[FFT.scala 53:18]
  wire [31:0] _GEN_880 = 8'h6f == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_879); // @[FFT.scala 53:18]
  wire [31:0] _GEN_881 = 8'h70 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_880); // @[FFT.scala 53:18]
  wire [31:0] _GEN_882 = 8'h71 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_881); // @[FFT.scala 53:18]
  wire [31:0] _GEN_883 = 8'h72 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_882); // @[FFT.scala 53:18]
  wire [31:0] _GEN_884 = 8'h73 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_883); // @[FFT.scala 53:18]
  wire [31:0] _GEN_885 = 8'h74 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_884); // @[FFT.scala 53:18]
  wire [31:0] _GEN_886 = 8'h75 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_885); // @[FFT.scala 53:18]
  wire [31:0] _GEN_887 = 8'h76 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_886); // @[FFT.scala 53:18]
  wire [31:0] _GEN_888 = 8'h77 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_887); // @[FFT.scala 53:18]
  wire [31:0] _GEN_889 = 8'h78 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_888); // @[FFT.scala 53:18]
  wire [31:0] _GEN_890 = 8'h79 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_889); // @[FFT.scala 53:18]
  wire [31:0] _GEN_891 = 8'h7a == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_890); // @[FFT.scala 53:18]
  wire [31:0] _GEN_892 = 8'h7b == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_891); // @[FFT.scala 53:18]
  wire [31:0] _GEN_893 = 8'h7c == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_892); // @[FFT.scala 53:18]
  wire [31:0] _GEN_894 = 8'h7d == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_893); // @[FFT.scala 53:18]
  wire [31:0] _GEN_895 = 8'h7e == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_894); // @[FFT.scala 53:18]
  wire [31:0] _GEN_896 = 8'h7f == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_895); // @[FFT.scala 53:18]
  wire [31:0] _GEN_897 = 8'h80 == cnt[7:0] ? $signed(-32'sh10000) : $signed(_GEN_896); // @[FFT.scala 53:18]
  wire [31:0] _GEN_898 = 8'h81 == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_897); // @[FFT.scala 53:18]
  wire [31:0] _GEN_899 = 8'h82 == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_898); // @[FFT.scala 53:18]
  wire [31:0] _GEN_900 = 8'h83 == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_899); // @[FFT.scala 53:18]
  wire [31:0] _GEN_901 = 8'h84 == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_900); // @[FFT.scala 53:18]
  wire [31:0] _GEN_902 = 8'h85 == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_901); // @[FFT.scala 53:18]
  wire [31:0] _GEN_903 = 8'h86 == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_902); // @[FFT.scala 53:18]
  wire [31:0] _GEN_904 = 8'h87 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_903); // @[FFT.scala 53:18]
  wire [31:0] _GEN_905 = 8'h88 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_904); // @[FFT.scala 53:18]
  wire [31:0] _GEN_906 = 8'h89 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_905); // @[FFT.scala 53:18]
  wire [31:0] _GEN_907 = 8'h8a == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_906); // @[FFT.scala 53:18]
  wire [31:0] _GEN_908 = 8'h8b == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_907); // @[FFT.scala 53:18]
  wire [31:0] _GEN_909 = 8'h8c == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_908); // @[FFT.scala 53:18]
  wire [31:0] _GEN_910 = 8'h8d == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_909); // @[FFT.scala 53:18]
  wire [31:0] _GEN_911 = 8'h8e == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_910); // @[FFT.scala 53:18]
  wire [31:0] _GEN_912 = 8'h8f == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_911); // @[FFT.scala 53:18]
  wire [31:0] _GEN_913 = 8'h90 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_912); // @[FFT.scala 53:18]
  wire [31:0] _GEN_914 = 8'h91 == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_913); // @[FFT.scala 53:18]
  wire [31:0] _GEN_915 = 8'h92 == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_914); // @[FFT.scala 53:18]
  wire [31:0] _GEN_916 = 8'h93 == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_915); // @[FFT.scala 53:18]
  wire [31:0] _GEN_917 = 8'h94 == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_916); // @[FFT.scala 53:18]
  wire [31:0] _GEN_918 = 8'h95 == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_917); // @[FFT.scala 53:18]
  wire [31:0] _GEN_919 = 8'h96 == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_918); // @[FFT.scala 53:18]
  wire [31:0] _GEN_920 = 8'h97 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_919); // @[FFT.scala 53:18]
  wire [31:0] _GEN_921 = 8'h98 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_920); // @[FFT.scala 53:18]
  wire [31:0] _GEN_922 = 8'h99 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_921); // @[FFT.scala 53:18]
  wire [31:0] _GEN_923 = 8'h9a == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_922); // @[FFT.scala 53:18]
  wire [31:0] _GEN_924 = 8'h9b == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_923); // @[FFT.scala 53:18]
  wire [31:0] _GEN_925 = 8'h9c == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_924); // @[FFT.scala 53:18]
  wire [31:0] _GEN_926 = 8'h9d == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_925); // @[FFT.scala 53:18]
  wire [31:0] _GEN_927 = 8'h9e == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_926); // @[FFT.scala 53:18]
  wire [31:0] _GEN_928 = 8'h9f == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_927); // @[FFT.scala 53:18]
  wire [31:0] _GEN_929 = 8'ha0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_928); // @[FFT.scala 53:18]
  wire [31:0] _GEN_930 = 8'ha1 == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_929); // @[FFT.scala 53:18]
  wire [31:0] _GEN_931 = 8'ha2 == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_930); // @[FFT.scala 53:18]
  wire [31:0] _GEN_932 = 8'ha3 == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_931); // @[FFT.scala 53:18]
  wire [31:0] _GEN_933 = 8'ha4 == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_932); // @[FFT.scala 53:18]
  wire [31:0] _GEN_934 = 8'ha5 == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_933); // @[FFT.scala 53:18]
  wire [31:0] _GEN_935 = 8'ha6 == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_934); // @[FFT.scala 53:18]
  wire [31:0] _GEN_936 = 8'ha7 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_935); // @[FFT.scala 53:18]
  wire [31:0] _GEN_937 = 8'ha8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_936); // @[FFT.scala 53:18]
  wire [31:0] _GEN_938 = 8'ha9 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_937); // @[FFT.scala 53:18]
  wire [31:0] _GEN_939 = 8'haa == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_938); // @[FFT.scala 53:18]
  wire [31:0] _GEN_940 = 8'hab == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_939); // @[FFT.scala 53:18]
  wire [31:0] _GEN_941 = 8'hac == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_940); // @[FFT.scala 53:18]
  wire [31:0] _GEN_942 = 8'had == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_941); // @[FFT.scala 53:18]
  wire [31:0] _GEN_943 = 8'hae == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_942); // @[FFT.scala 53:18]
  wire [31:0] _GEN_944 = 8'haf == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_943); // @[FFT.scala 53:18]
  wire [31:0] _GEN_945 = 8'hb0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_944); // @[FFT.scala 53:18]
  wire [31:0] _GEN_946 = 8'hb1 == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_945); // @[FFT.scala 53:18]
  wire [31:0] _GEN_947 = 8'hb2 == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_946); // @[FFT.scala 53:18]
  wire [31:0] _GEN_948 = 8'hb3 == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_947); // @[FFT.scala 53:18]
  wire [31:0] _GEN_949 = 8'hb4 == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_948); // @[FFT.scala 53:18]
  wire [31:0] _GEN_950 = 8'hb5 == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_949); // @[FFT.scala 53:18]
  wire [31:0] _GEN_951 = 8'hb6 == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_950); // @[FFT.scala 53:18]
  wire [31:0] _GEN_952 = 8'hb7 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_951); // @[FFT.scala 53:18]
  wire [31:0] _GEN_953 = 8'hb8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_952); // @[FFT.scala 53:18]
  wire [31:0] _GEN_954 = 8'hb9 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_953); // @[FFT.scala 53:18]
  wire [31:0] _GEN_955 = 8'hba == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_954); // @[FFT.scala 53:18]
  wire [31:0] _GEN_956 = 8'hbb == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_955); // @[FFT.scala 53:18]
  wire [31:0] _GEN_957 = 8'hbc == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_956); // @[FFT.scala 53:18]
  wire [31:0] _GEN_958 = 8'hbd == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_957); // @[FFT.scala 53:18]
  wire [31:0] _GEN_959 = 8'hbe == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_958); // @[FFT.scala 53:18]
  wire [31:0] _GEN_960 = 8'hbf == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_959); // @[FFT.scala 53:18]
  wire [31:0] _GEN_961 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_960); // @[FFT.scala 53:18]
  wire [31:0] _GEN_962 = 8'hc1 == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_961); // @[FFT.scala 53:18]
  wire [31:0] _GEN_963 = 8'hc2 == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_962); // @[FFT.scala 53:18]
  wire [31:0] _GEN_964 = 8'hc3 == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_963); // @[FFT.scala 53:18]
  wire [31:0] _GEN_965 = 8'hc4 == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_964); // @[FFT.scala 53:18]
  wire [31:0] _GEN_966 = 8'hc5 == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_965); // @[FFT.scala 53:18]
  wire [31:0] _GEN_967 = 8'hc6 == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_966); // @[FFT.scala 53:18]
  wire [31:0] _GEN_968 = 8'hc7 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_967); // @[FFT.scala 53:18]
  wire [31:0] _GEN_969 = 8'hc8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_968); // @[FFT.scala 53:18]
  wire [31:0] _GEN_970 = 8'hc9 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_969); // @[FFT.scala 53:18]
  wire [31:0] _GEN_971 = 8'hca == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_970); // @[FFT.scala 53:18]
  wire [31:0] _GEN_972 = 8'hcb == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_971); // @[FFT.scala 53:18]
  wire [31:0] _GEN_973 = 8'hcc == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_972); // @[FFT.scala 53:18]
  wire [31:0] _GEN_974 = 8'hcd == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_973); // @[FFT.scala 53:18]
  wire [31:0] _GEN_975 = 8'hce == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_974); // @[FFT.scala 53:18]
  wire [31:0] _GEN_976 = 8'hcf == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_975); // @[FFT.scala 53:18]
  wire [31:0] _GEN_977 = 8'hd0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_976); // @[FFT.scala 53:18]
  wire [31:0] _GEN_978 = 8'hd1 == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_977); // @[FFT.scala 53:18]
  wire [31:0] _GEN_979 = 8'hd2 == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_978); // @[FFT.scala 53:18]
  wire [31:0] _GEN_980 = 8'hd3 == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_979); // @[FFT.scala 53:18]
  wire [31:0] _GEN_981 = 8'hd4 == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_980); // @[FFT.scala 53:18]
  wire [31:0] _GEN_982 = 8'hd5 == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_981); // @[FFT.scala 53:18]
  wire [31:0] _GEN_983 = 8'hd6 == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_982); // @[FFT.scala 53:18]
  wire [31:0] _GEN_984 = 8'hd7 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_983); // @[FFT.scala 53:18]
  wire [31:0] _GEN_985 = 8'hd8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_984); // @[FFT.scala 53:18]
  wire [31:0] _GEN_986 = 8'hd9 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_985); // @[FFT.scala 53:18]
  wire [31:0] _GEN_987 = 8'hda == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_986); // @[FFT.scala 53:18]
  wire [31:0] _GEN_988 = 8'hdb == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_987); // @[FFT.scala 53:18]
  wire [31:0] _GEN_989 = 8'hdc == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_988); // @[FFT.scala 53:18]
  wire [31:0] _GEN_990 = 8'hdd == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_989); // @[FFT.scala 53:18]
  wire [31:0] _GEN_991 = 8'hde == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_990); // @[FFT.scala 53:18]
  wire [31:0] _GEN_992 = 8'hdf == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_991); // @[FFT.scala 53:18]
  wire [31:0] _GEN_993 = 8'he0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_992); // @[FFT.scala 53:18]
  wire [31:0] _GEN_994 = 8'he1 == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_993); // @[FFT.scala 53:18]
  wire [31:0] _GEN_995 = 8'he2 == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_994); // @[FFT.scala 53:18]
  wire [31:0] _GEN_996 = 8'he3 == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_995); // @[FFT.scala 53:18]
  wire [31:0] _GEN_997 = 8'he4 == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_996); // @[FFT.scala 53:18]
  wire [31:0] _GEN_998 = 8'he5 == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_997); // @[FFT.scala 53:18]
  wire [31:0] _GEN_999 = 8'he6 == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_998); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1000 = 8'he7 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_999); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1001 = 8'he8 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_1000); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1002 = 8'he9 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_1001); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1003 = 8'hea == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_1002); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1004 = 8'heb == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_1003); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1005 = 8'hec == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_1004); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1006 = 8'hed == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_1005); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1007 = 8'hee == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_1006); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1008 = 8'hef == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_1007); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1009 = 8'hf0 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_1008); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1010 = 8'hf1 == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_1009); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1011 = 8'hf2 == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1010); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1012 = 8'hf3 == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_1011); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1013 = 8'hf4 == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_1012); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1014 = 8'hf5 == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_1013); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1015 = 8'hf6 == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_1014); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1016 = 8'hf7 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_1015); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1017 = 8'hf8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_1016); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1018 = 8'hf9 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_1017); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1019 = 8'hfa == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_1018); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1020 = 8'hfb == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_1019); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1021 = 8'hfc == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_1020); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1022 = 8'hfd == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_1021); // @[FFT.scala 53:18]
  wire [31:0] _GEN_1023 = 8'hfe == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_1022); // @[FFT.scala 53:18]
  reg [31:0] _T_153_re; // @[Reg.scala 15:16]
  reg [31:0] _T_154_re; // @[Reg.scala 15:16]
  reg [31:0] _T_155_re; // @[Reg.scala 15:16]
  reg [31:0] _T_156_re; // @[Reg.scala 15:16]
  reg [31:0] _T_157_re; // @[Reg.scala 15:16]
  reg [31:0] _T_158_re; // @[Reg.scala 15:16]
  reg [31:0] _T_159_re; // @[Reg.scala 15:16]
  reg [31:0] _T_160_re; // @[Reg.scala 15:16]
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _T_533_re; // @[Reg.scala 15:16]
  reg [31:0] _T_533_im; // @[Reg.scala 15:16]
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _T_536_re; // @[Reg.scala 15:16]
  reg [31:0] _T_536_im; // @[Reg.scala 15:16]
  reg [31:0] _T_537_re; // @[Reg.scala 15:16]
  reg [31:0] _T_537_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_1794 = 7'h1 == cnt[6:0] ? $signed(32'shffec) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1795 = 7'h2 == cnt[6:0] ? $signed(32'shffb1) : $signed(_GEN_1794); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1796 = 7'h3 == cnt[6:0] ? $signed(32'shff4e) : $signed(_GEN_1795); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1797 = 7'h4 == cnt[6:0] ? $signed(32'shfec4) : $signed(_GEN_1796); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1798 = 7'h5 == cnt[6:0] ? $signed(32'shfe13) : $signed(_GEN_1797); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1799 = 7'h6 == cnt[6:0] ? $signed(32'shfd3b) : $signed(_GEN_1798); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1800 = 7'h7 == cnt[6:0] ? $signed(32'shfc3b) : $signed(_GEN_1799); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1801 = 7'h8 == cnt[6:0] ? $signed(32'shfb15) : $signed(_GEN_1800); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1802 = 7'h9 == cnt[6:0] ? $signed(32'shf9c8) : $signed(_GEN_1801); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1803 = 7'ha == cnt[6:0] ? $signed(32'shf854) : $signed(_GEN_1802); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1804 = 7'hb == cnt[6:0] ? $signed(32'shf6ba) : $signed(_GEN_1803); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1805 = 7'hc == cnt[6:0] ? $signed(32'shf4fa) : $signed(_GEN_1804); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1806 = 7'hd == cnt[6:0] ? $signed(32'shf314) : $signed(_GEN_1805); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1807 = 7'he == cnt[6:0] ? $signed(32'shf109) : $signed(_GEN_1806); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1808 = 7'hf == cnt[6:0] ? $signed(32'sheed9) : $signed(_GEN_1807); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1809 = 7'h10 == cnt[6:0] ? $signed(32'shec83) : $signed(_GEN_1808); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1810 = 7'h11 == cnt[6:0] ? $signed(32'shea0a) : $signed(_GEN_1809); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1811 = 7'h12 == cnt[6:0] ? $signed(32'she76c) : $signed(_GEN_1810); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1812 = 7'h13 == cnt[6:0] ? $signed(32'she4aa) : $signed(_GEN_1811); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1813 = 7'h14 == cnt[6:0] ? $signed(32'she1c6) : $signed(_GEN_1812); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1814 = 7'h15 == cnt[6:0] ? $signed(32'shdebe) : $signed(_GEN_1813); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1815 = 7'h16 == cnt[6:0] ? $signed(32'shdb94) : $signed(_GEN_1814); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1816 = 7'h17 == cnt[6:0] ? $signed(32'shd848) : $signed(_GEN_1815); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1817 = 7'h18 == cnt[6:0] ? $signed(32'shd4db) : $signed(_GEN_1816); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1818 = 7'h19 == cnt[6:0] ? $signed(32'shd14d) : $signed(_GEN_1817); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1819 = 7'h1a == cnt[6:0] ? $signed(32'shcd9f) : $signed(_GEN_1818); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1820 = 7'h1b == cnt[6:0] ? $signed(32'shc9d1) : $signed(_GEN_1819); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1821 = 7'h1c == cnt[6:0] ? $signed(32'shc5e4) : $signed(_GEN_1820); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1822 = 7'h1d == cnt[6:0] ? $signed(32'shc1d8) : $signed(_GEN_1821); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1823 = 7'h1e == cnt[6:0] ? $signed(32'shbdaf) : $signed(_GEN_1822); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1824 = 7'h1f == cnt[6:0] ? $signed(32'shb968) : $signed(_GEN_1823); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1825 = 7'h20 == cnt[6:0] ? $signed(32'shb505) : $signed(_GEN_1824); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1826 = 7'h21 == cnt[6:0] ? $signed(32'shb086) : $signed(_GEN_1825); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1827 = 7'h22 == cnt[6:0] ? $signed(32'shabeb) : $signed(_GEN_1826); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1828 = 7'h23 == cnt[6:0] ? $signed(32'sha736) : $signed(_GEN_1827); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1829 = 7'h24 == cnt[6:0] ? $signed(32'sha268) : $signed(_GEN_1828); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1830 = 7'h25 == cnt[6:0] ? $signed(32'sh9d80) : $signed(_GEN_1829); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1831 = 7'h26 == cnt[6:0] ? $signed(32'sh9880) : $signed(_GEN_1830); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1832 = 7'h27 == cnt[6:0] ? $signed(32'sh9368) : $signed(_GEN_1831); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1833 = 7'h28 == cnt[6:0] ? $signed(32'sh8e3a) : $signed(_GEN_1832); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1834 = 7'h29 == cnt[6:0] ? $signed(32'sh88f6) : $signed(_GEN_1833); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1835 = 7'h2a == cnt[6:0] ? $signed(32'sh839c) : $signed(_GEN_1834); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1836 = 7'h2b == cnt[6:0] ? $signed(32'sh7e2f) : $signed(_GEN_1835); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1837 = 7'h2c == cnt[6:0] ? $signed(32'sh78ad) : $signed(_GEN_1836); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1838 = 7'h2d == cnt[6:0] ? $signed(32'sh731a) : $signed(_GEN_1837); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1839 = 7'h2e == cnt[6:0] ? $signed(32'sh6d74) : $signed(_GEN_1838); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1840 = 7'h2f == cnt[6:0] ? $signed(32'sh67be) : $signed(_GEN_1839); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1841 = 7'h30 == cnt[6:0] ? $signed(32'sh61f8) : $signed(_GEN_1840); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1842 = 7'h31 == cnt[6:0] ? $signed(32'sh5c22) : $signed(_GEN_1841); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1843 = 7'h32 == cnt[6:0] ? $signed(32'sh563e) : $signed(_GEN_1842); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1844 = 7'h33 == cnt[6:0] ? $signed(32'sh504d) : $signed(_GEN_1843); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1845 = 7'h34 == cnt[6:0] ? $signed(32'sh4a50) : $signed(_GEN_1844); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1846 = 7'h35 == cnt[6:0] ? $signed(32'sh4447) : $signed(_GEN_1845); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1847 = 7'h36 == cnt[6:0] ? $signed(32'sh3e34) : $signed(_GEN_1846); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1848 = 7'h37 == cnt[6:0] ? $signed(32'sh3817) : $signed(_GEN_1847); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1849 = 7'h38 == cnt[6:0] ? $signed(32'sh31f1) : $signed(_GEN_1848); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1850 = 7'h39 == cnt[6:0] ? $signed(32'sh2bc4) : $signed(_GEN_1849); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1851 = 7'h3a == cnt[6:0] ? $signed(32'sh2590) : $signed(_GEN_1850); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1852 = 7'h3b == cnt[6:0] ? $signed(32'sh1f56) : $signed(_GEN_1851); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1853 = 7'h3c == cnt[6:0] ? $signed(32'sh1918) : $signed(_GEN_1852); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1854 = 7'h3d == cnt[6:0] ? $signed(32'sh12d5) : $signed(_GEN_1853); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1855 = 7'h3e == cnt[6:0] ? $signed(32'shc90) : $signed(_GEN_1854); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1856 = 7'h3f == cnt[6:0] ? $signed(32'sh648) : $signed(_GEN_1855); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1857 = 7'h40 == cnt[6:0] ? $signed(32'sh0) : $signed(_GEN_1856); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1858 = 7'h41 == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_1857); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1859 = 7'h42 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_1858); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1860 = 7'h43 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_1859); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1861 = 7'h44 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_1860); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1862 = 7'h45 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_1861); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1863 = 7'h46 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_1862); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1864 = 7'h47 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1863); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1865 = 7'h48 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_1864); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1866 = 7'h49 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_1865); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1867 = 7'h4a == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_1866); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1868 = 7'h4b == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_1867); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1869 = 7'h4c == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_1868); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1870 = 7'h4d == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_1869); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1871 = 7'h4e == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_1870); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1872 = 7'h4f == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_1871); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1873 = 7'h50 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_1872); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1874 = 7'h51 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_1873); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1875 = 7'h52 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_1874); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1876 = 7'h53 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_1875); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1877 = 7'h54 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_1876); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1878 = 7'h55 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_1877); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1879 = 7'h56 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_1878); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1880 = 7'h57 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_1879); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1881 = 7'h58 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1880); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1882 = 7'h59 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_1881); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1883 = 7'h5a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_1882); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1884 = 7'h5b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_1883); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1885 = 7'h5c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_1884); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1886 = 7'h5d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_1885); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1887 = 7'h5e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_1886); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1888 = 7'h5f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_1887); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1889 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_1888); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1890 = 7'h61 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_1889); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1891 = 7'h62 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_1890); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1892 = 7'h63 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_1891); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1893 = 7'h64 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_1892); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1894 = 7'h65 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_1893); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1895 = 7'h66 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_1894); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1896 = 7'h67 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_1895); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1897 = 7'h68 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_1896); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1898 = 7'h69 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_1897); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1899 = 7'h6a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_1898); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1900 = 7'h6b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_1899); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1901 = 7'h6c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_1900); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1902 = 7'h6d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_1901); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1903 = 7'h6e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_1902); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1904 = 7'h6f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_1903); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1905 = 7'h70 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_1904); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1906 = 7'h71 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_1905); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1907 = 7'h72 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_1906); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1908 = 7'h73 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_1907); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1909 = 7'h74 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_1908); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1910 = 7'h75 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_1909); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1911 = 7'h76 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_1910); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1912 = 7'h77 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_1911); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1913 = 7'h78 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_1912); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1914 = 7'h79 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_1913); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1915 = 7'h7a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_1914); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1916 = 7'h7b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_1915); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1917 = 7'h7c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_1916); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1918 = 7'h7d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_1917); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1919 = 7'h7e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_1918); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2178 = 7'h1 == cnt[6:0] ? $signed(-32'sh648) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2179 = 7'h2 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_2178); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2180 = 7'h3 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_2179); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2181 = 7'h4 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_2180); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2182 = 7'h5 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_2181); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2183 = 7'h6 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_2182); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2184 = 7'h7 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2183); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2185 = 7'h8 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_2184); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2186 = 7'h9 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_2185); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2187 = 7'ha == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_2186); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2188 = 7'hb == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_2187); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2189 = 7'hc == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_2188); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2190 = 7'hd == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_2189); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2191 = 7'he == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_2190); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2192 = 7'hf == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_2191); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2193 = 7'h10 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_2192); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2194 = 7'h11 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_2193); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2195 = 7'h12 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_2194); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2196 = 7'h13 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_2195); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2197 = 7'h14 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_2196); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2198 = 7'h15 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2197); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2199 = 7'h16 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_2198); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2200 = 7'h17 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_2199); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2201 = 7'h18 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2200); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2202 = 7'h19 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_2201); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2203 = 7'h1a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_2202); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2204 = 7'h1b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_2203); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2205 = 7'h1c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_2204); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2206 = 7'h1d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_2205); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2207 = 7'h1e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_2206); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2208 = 7'h1f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_2207); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2209 = 7'h20 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_2208); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2210 = 7'h21 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_2209); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2211 = 7'h22 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_2210); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2212 = 7'h23 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_2211); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2213 = 7'h24 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_2212); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2214 = 7'h25 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_2213); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2215 = 7'h26 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_2214); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2216 = 7'h27 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_2215); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2217 = 7'h28 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_2216); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2218 = 7'h29 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_2217); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2219 = 7'h2a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_2218); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2220 = 7'h2b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_2219); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2221 = 7'h2c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_2220); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2222 = 7'h2d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_2221); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2223 = 7'h2e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_2222); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2224 = 7'h2f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_2223); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2225 = 7'h30 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_2224); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2226 = 7'h31 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_2225); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2227 = 7'h32 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_2226); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2228 = 7'h33 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_2227); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2229 = 7'h34 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_2228); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2230 = 7'h35 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_2229); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2231 = 7'h36 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_2230); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2232 = 7'h37 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_2231); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2233 = 7'h38 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_2232); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2234 = 7'h39 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_2233); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2235 = 7'h3a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_2234); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2236 = 7'h3b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_2235); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2237 = 7'h3c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_2236); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2238 = 7'h3d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_2237); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2239 = 7'h3e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_2238); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2240 = 7'h3f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_2239); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2241 = 7'h40 == cnt[6:0] ? $signed(-32'sh10000) : $signed(_GEN_2240); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2242 = 7'h41 == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_2241); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2243 = 7'h42 == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_2242); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2244 = 7'h43 == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_2243); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2245 = 7'h44 == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_2244); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2246 = 7'h45 == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_2245); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2247 = 7'h46 == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_2246); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2248 = 7'h47 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_2247); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2249 = 7'h48 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_2248); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2250 = 7'h49 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_2249); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2251 = 7'h4a == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_2250); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2252 = 7'h4b == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_2251); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2253 = 7'h4c == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_2252); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2254 = 7'h4d == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_2253); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2255 = 7'h4e == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_2254); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2256 = 7'h4f == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_2255); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2257 = 7'h50 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_2256); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2258 = 7'h51 == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_2257); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2259 = 7'h52 == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_2258); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2260 = 7'h53 == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_2259); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2261 = 7'h54 == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_2260); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2262 = 7'h55 == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_2261); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2263 = 7'h56 == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_2262); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2264 = 7'h57 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_2263); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2265 = 7'h58 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_2264); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2266 = 7'h59 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_2265); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2267 = 7'h5a == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_2266); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2268 = 7'h5b == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_2267); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2269 = 7'h5c == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_2268); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2270 = 7'h5d == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_2269); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2271 = 7'h5e == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_2270); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2272 = 7'h5f == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_2271); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2273 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_2272); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2274 = 7'h61 == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_2273); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2275 = 7'h62 == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_2274); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2276 = 7'h63 == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_2275); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2277 = 7'h64 == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_2276); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2278 = 7'h65 == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_2277); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2279 = 7'h66 == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_2278); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2280 = 7'h67 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_2279); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2281 = 7'h68 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2280); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2282 = 7'h69 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_2281); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2283 = 7'h6a == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_2282); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2284 = 7'h6b == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2283); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2285 = 7'h6c == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_2284); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2286 = 7'h6d == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_2285); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2287 = 7'h6e == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_2286); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2288 = 7'h6f == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_2287); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2289 = 7'h70 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_2288); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2290 = 7'h71 == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_2289); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2291 = 7'h72 == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_2290); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2292 = 7'h73 == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_2291); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2293 = 7'h74 == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_2292); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2294 = 7'h75 == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_2293); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2295 = 7'h76 == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_2294); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2296 = 7'h77 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_2295); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2297 = 7'h78 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_2296); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2298 = 7'h79 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2297); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2299 = 7'h7a == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_2298); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2300 = 7'h7b == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_2299); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2301 = 7'h7c == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_2300); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2302 = 7'h7d == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_2301); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2303 = 7'h7e == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_2302); // @[FFT.scala 53:18]
  reg [31:0] _T_546_re; // @[Reg.scala 15:16]
  reg [31:0] _T_546_im; // @[Reg.scala 15:16]
  reg [31:0] _T_547_re; // @[Reg.scala 15:16]
  reg [31:0] _T_547_im; // @[Reg.scala 15:16]
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _T_663_re; // @[Reg.scala 15:16]
  reg [31:0] _T_663_im; // @[Reg.scala 15:16]
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _T_671_re; // @[Reg.scala 15:16]
  reg [31:0] _T_671_im; // @[Reg.scala 15:16]
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _T_673_re; // @[Reg.scala 15:16]
  reg [31:0] _T_673_im; // @[Reg.scala 15:16]
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _T_676_re; // @[Reg.scala 15:16]
  reg [31:0] _T_676_im; // @[Reg.scala 15:16]
  reg [31:0] _T_677_re; // @[Reg.scala 15:16]
  reg [31:0] _T_677_im; // @[Reg.scala 15:16]
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _T_728_re; // @[Reg.scala 15:16]
  reg [31:0] _T_728_im; // @[Reg.scala 15:16]
  reg [31:0] _T_729_re; // @[Reg.scala 15:16]
  reg [31:0] _T_729_im; // @[Reg.scala 15:16]
  reg [31:0] _T_730_re; // @[Reg.scala 15:16]
  reg [31:0] _T_730_im; // @[Reg.scala 15:16]
  reg [31:0] _T_731_re; // @[Reg.scala 15:16]
  reg [31:0] _T_731_im; // @[Reg.scala 15:16]
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  reg [31:0] _T_736_re; // @[Reg.scala 15:16]
  reg [31:0] _T_736_im; // @[Reg.scala 15:16]
  reg [31:0] _T_737_re; // @[Reg.scala 15:16]
  reg [31:0] _T_737_im; // @[Reg.scala 15:16]
  reg [31:0] _T_738_re; // @[Reg.scala 15:16]
  reg [31:0] _T_738_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_2690 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2691 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_2690); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2692 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_2691); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2693 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_2692); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2694 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_2693); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2695 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_2694); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2696 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_2695); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2697 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_2696); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2698 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_2697); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2699 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_2698); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2700 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_2699); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2701 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_2700); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2702 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_2701); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2703 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_2702); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2704 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_2703); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2705 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_2704); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2706 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_2705); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2707 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_2706); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2708 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_2707); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2709 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_2708); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2710 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_2709); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2711 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_2710); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2712 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_2711); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2713 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_2712); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2714 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_2713); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2715 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_2714); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2716 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_2715); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2717 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_2716); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2718 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_2717); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2719 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_2718); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2720 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_2719); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2721 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_2720); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2722 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_2721); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2723 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2722); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2724 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2723); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2725 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2724); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2726 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2725); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2727 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2726); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2728 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2727); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2729 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2728); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2730 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2729); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2731 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2730); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2732 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2731); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2733 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2732); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2734 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2733); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2735 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2734); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2736 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2735); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2737 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2736); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2738 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2737); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2739 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2738); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2740 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2739); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2741 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2740); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2742 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2741); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2743 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2742); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2744 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2743); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2745 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2744); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2746 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2745); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2747 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2746); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2748 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2747); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2749 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2748); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2750 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2749); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2751 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2750); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2882 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2883 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2882); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2884 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2883); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2885 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2884); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2886 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2885); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2887 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2886); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2888 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2887); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2889 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2888); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2890 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2889); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2891 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2890); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2892 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2891); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2893 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2892); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2894 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2893); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2895 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2894); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2896 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2895); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2897 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2896); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2898 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2897); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2899 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2898); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2900 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2899); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2901 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2900); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2902 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2901); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2903 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2902); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2904 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2903); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2905 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2904); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2906 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2905); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2907 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2906); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2908 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2907); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2909 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2908); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2910 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2909); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2911 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2910); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2912 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2911); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2913 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_2912); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2914 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2913); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2915 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2914); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2916 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2915); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2917 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2916); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2918 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2917); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2919 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2918); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2920 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2919); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2921 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2920); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2922 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2921); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2923 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2922); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2924 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2923); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2925 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2924); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2926 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2925); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2927 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2926); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2928 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2927); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2929 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2928); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2930 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2929); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2931 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2930); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2932 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2931); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2933 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2932); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2934 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2933); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2935 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2934); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2936 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2935); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2937 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2936); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2938 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2937); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2939 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2938); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2940 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2939); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2941 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2940); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2942 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2941); // @[FFT.scala 53:18]
  wire [31:0] _GEN_2943 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2942); // @[FFT.scala 53:18]
  reg [31:0] _T_747_re; // @[Reg.scala 15:16]
  reg [31:0] _T_747_im; // @[Reg.scala 15:16]
  reg [31:0] _T_748_re; // @[Reg.scala 15:16]
  reg [31:0] _T_748_im; // @[Reg.scala 15:16]
  reg [31:0] _T_749_re; // @[Reg.scala 15:16]
  reg [31:0] _T_749_im; // @[Reg.scala 15:16]
  reg [31:0] _T_750_re; // @[Reg.scala 15:16]
  reg [31:0] _T_750_im; // @[Reg.scala 15:16]
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _T_796_re; // @[Reg.scala 15:16]
  reg [31:0] _T_796_im; // @[Reg.scala 15:16]
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _T_808_re; // @[Reg.scala 15:16]
  reg [31:0] _T_808_im; // @[Reg.scala 15:16]
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _T_815_re; // @[Reg.scala 15:16]
  reg [31:0] _T_815_im; // @[Reg.scala 15:16]
  reg [31:0] _T_816_re; // @[Reg.scala 15:16]
  reg [31:0] _T_816_im; // @[Reg.scala 15:16]
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _T_829_re; // @[Reg.scala 15:16]
  reg [31:0] _T_829_im; // @[Reg.scala 15:16]
  reg [31:0] _T_830_re; // @[Reg.scala 15:16]
  reg [31:0] _T_830_im; // @[Reg.scala 15:16]
  reg [31:0] _T_831_re; // @[Reg.scala 15:16]
  reg [31:0] _T_831_im; // @[Reg.scala 15:16]
  reg [31:0] _T_832_re; // @[Reg.scala 15:16]
  reg [31:0] _T_832_im; // @[Reg.scala 15:16]
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  reg [31:0] _T_841_re; // @[Reg.scala 15:16]
  reg [31:0] _T_841_im; // @[Reg.scala 15:16]
  reg [31:0] _T_842_re; // @[Reg.scala 15:16]
  reg [31:0] _T_842_im; // @[Reg.scala 15:16]
  reg [31:0] _T_843_re; // @[Reg.scala 15:16]
  reg [31:0] _T_843_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3138 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3139 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_3138); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3140 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_3139); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3141 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_3140); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3142 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_3141); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3143 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_3142); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3144 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_3143); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3145 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_3144); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3146 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_3145); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3147 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_3146); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3148 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_3147); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3149 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_3148); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3150 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_3149); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3151 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_3150); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3152 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_3151); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3153 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_3152); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3154 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_3153); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3155 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_3154); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3156 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_3155); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3157 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_3156); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3158 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_3157); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3159 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3158); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3160 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_3159); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3161 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_3160); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3162 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_3161); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3163 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_3162); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3164 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_3163); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3165 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_3164); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3166 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_3165); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3167 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_3166); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3234 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3235 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_3234); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3236 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_3235); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3237 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_3236); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3238 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_3237); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3239 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3238); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3240 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_3239); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3241 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_3240); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3242 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_3241); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3243 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_3242); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3244 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_3243); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3245 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_3244); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3246 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_3245); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3247 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_3246); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3248 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_3247); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3249 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_3248); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3250 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_3249); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3251 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_3250); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3252 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_3251); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3253 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_3252); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3254 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_3253); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3255 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_3254); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3256 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_3255); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3257 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_3256); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3258 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_3257); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3259 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3258); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3260 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_3259); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3261 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_3260); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3262 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_3261); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3263 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_3262); // @[FFT.scala 53:18]
  reg [31:0] _T_852_re; // @[Reg.scala 15:16]
  reg [31:0] _T_852_im; // @[Reg.scala 15:16]
  reg [31:0] _T_853_re; // @[Reg.scala 15:16]
  reg [31:0] _T_853_im; // @[Reg.scala 15:16]
  reg [31:0] _T_854_re; // @[Reg.scala 15:16]
  reg [31:0] _T_854_im; // @[Reg.scala 15:16]
  reg [31:0] _T_855_re; // @[Reg.scala 15:16]
  reg [31:0] _T_855_im; // @[Reg.scala 15:16]
  reg [31:0] _T_856_re; // @[Reg.scala 15:16]
  reg [31:0] _T_856_im; // @[Reg.scala 15:16]
  reg [31:0] _T_857_re; // @[Reg.scala 15:16]
  reg [31:0] _T_857_im; // @[Reg.scala 15:16]
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _T_865_re; // @[Reg.scala 15:16]
  reg [31:0] _T_865_im; // @[Reg.scala 15:16]
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _T_881_re; // @[Reg.scala 15:16]
  reg [31:0] _T_881_im; // @[Reg.scala 15:16]
  reg [31:0] _T_882_re; // @[Reg.scala 15:16]
  reg [31:0] _T_882_im; // @[Reg.scala 15:16]
  reg [31:0] _T_883_re; // @[Reg.scala 15:16]
  reg [31:0] _T_883_im; // @[Reg.scala 15:16]
  reg [31:0] _T_885_re; // @[Reg.scala 15:16]
  reg [31:0] _T_885_im; // @[Reg.scala 15:16]
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _T_890_re; // @[Reg.scala 15:16]
  reg [31:0] _T_890_im; // @[Reg.scala 15:16]
  reg [31:0] _T_891_re; // @[Reg.scala 15:16]
  reg [31:0] _T_891_im; // @[Reg.scala 15:16]
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  reg [31:0] _T_898_re; // @[Reg.scala 15:16]
  reg [31:0] _T_898_im; // @[Reg.scala 15:16]
  reg [31:0] _T_899_re; // @[Reg.scala 15:16]
  reg [31:0] _T_899_im; // @[Reg.scala 15:16]
  reg [31:0] _T_900_re; // @[Reg.scala 15:16]
  reg [31:0] _T_900_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3362 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3363 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_3362); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3364 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_3363); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3365 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_3364); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3366 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_3365); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3367 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_3366); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3368 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_3367); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3369 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_3368); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3370 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_3369); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3371 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_3370); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3372 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3371); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3373 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_3372); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3374 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_3373); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3375 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_3374); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3410 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3411 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_3410); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3412 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3411); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3413 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_3412); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3414 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_3413); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3415 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_3414); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3416 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_3415); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3417 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_3416); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3418 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_3417); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3419 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_3418); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3420 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_3419); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3421 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_3420); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3422 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3421); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3423 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_3422); // @[FFT.scala 53:18]
  reg [31:0] _T_909_re; // @[Reg.scala 15:16]
  reg [31:0] _T_909_im; // @[Reg.scala 15:16]
  reg [31:0] _T_910_re; // @[Reg.scala 15:16]
  reg [31:0] _T_910_im; // @[Reg.scala 15:16]
  reg [31:0] _T_911_re; // @[Reg.scala 15:16]
  reg [31:0] _T_911_im; // @[Reg.scala 15:16]
  reg [31:0] _T_912_re; // @[Reg.scala 15:16]
  reg [31:0] _T_912_im; // @[Reg.scala 15:16]
  reg [31:0] _T_913_re; // @[Reg.scala 15:16]
  reg [31:0] _T_913_im; // @[Reg.scala 15:16]
  reg [31:0] _T_914_re; // @[Reg.scala 15:16]
  reg [31:0] _T_914_im; // @[Reg.scala 15:16]
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _T_922_re; // @[Reg.scala 15:16]
  reg [31:0] _T_922_im; // @[Reg.scala 15:16]
  reg [31:0] _T_923_re; // @[Reg.scala 15:16]
  reg [31:0] _T_923_im; // @[Reg.scala 15:16]
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _T_928_re; // @[Reg.scala 15:16]
  reg [31:0] _T_928_im; // @[Reg.scala 15:16]
  reg [31:0] _T_929_re; // @[Reg.scala 15:16]
  reg [31:0] _T_929_im; // @[Reg.scala 15:16]
  reg [31:0] _T_930_re; // @[Reg.scala 15:16]
  reg [31:0] _T_930_im; // @[Reg.scala 15:16]
  reg [31:0] _T_931_re; // @[Reg.scala 15:16]
  reg [31:0] _T_931_im; // @[Reg.scala 15:16]
  reg [31:0] _T_932_re; // @[Reg.scala 15:16]
  reg [31:0] _T_932_im; // @[Reg.scala 15:16]
  reg [31:0] _T_933_re; // @[Reg.scala 15:16]
  reg [31:0] _T_933_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3474 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3475 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_3474); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3476 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_3475); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3477 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_3476); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3478 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_3477); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3479 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_3478); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3498 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3499 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_3498); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3500 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_3499); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3501 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_3500); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3502 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_3501); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3503 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_3502); // @[FFT.scala 53:18]
  reg [31:0] _T_942_re; // @[Reg.scala 15:16]
  reg [31:0] _T_942_im; // @[Reg.scala 15:16]
  reg [31:0] _T_943_re; // @[Reg.scala 15:16]
  reg [31:0] _T_943_im; // @[Reg.scala 15:16]
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _T_945_re; // @[Reg.scala 15:16]
  reg [31:0] _T_945_im; // @[Reg.scala 15:16]
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _T_947_re; // @[Reg.scala 15:16]
  reg [31:0] _T_947_im; // @[Reg.scala 15:16]
  reg [31:0] _T_948_re; // @[Reg.scala 15:16]
  reg [31:0] _T_948_im; // @[Reg.scala 15:16]
  reg [31:0] _T_949_re; // @[Reg.scala 15:16]
  reg [31:0] _T_949_im; // @[Reg.scala 15:16]
  reg [31:0] _T_951_re; // @[Reg.scala 15:16]
  reg [31:0] _T_951_im; // @[Reg.scala 15:16]
  reg [31:0] _T_952_re; // @[Reg.scala 15:16]
  reg [31:0] _T_952_im; // @[Reg.scala 15:16]
  reg [31:0] _T_953_re; // @[Reg.scala 15:16]
  reg [31:0] _T_953_im; // @[Reg.scala 15:16]
  reg [31:0] _T_954_re; // @[Reg.scala 15:16]
  reg [31:0] _T_954_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3530 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3531 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_3530); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3542 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 53:18]
  wire [31:0] _GEN_3543 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_3542); // @[FFT.scala 53:18]
  reg [31:0] _T_963_re; // @[Reg.scala 15:16]
  reg [31:0] _T_963_im; // @[Reg.scala 15:16]
  reg [31:0] _T_964_re; // @[Reg.scala 15:16]
  reg [31:0] _T_964_im; // @[Reg.scala 15:16]
  reg [31:0] _T_965_re; // @[Reg.scala 15:16]
  reg [31:0] _T_965_im; // @[Reg.scala 15:16]
  reg [31:0] _T_966_re; // @[Reg.scala 15:16]
  reg [31:0] _T_966_im; // @[Reg.scala 15:16]
  reg [31:0] _T_968_re; // @[Reg.scala 15:16]
  reg [31:0] _T_968_im; // @[Reg.scala 15:16]
  reg [31:0] _T_969_re; // @[Reg.scala 15:16]
  reg [31:0] _T_969_im; // @[Reg.scala 15:16]
  reg [31:0] _T_978_re; // @[Reg.scala 15:16]
  reg [31:0] _T_978_im; // @[Reg.scala 15:16]
  reg [31:0] _T_979_re; // @[Reg.scala 15:16]
  reg [31:0] _T_979_im; // @[Reg.scala 15:16]
  reg [31:0] _T_981_re; // @[Reg.scala 15:16]
  reg [31:0] _T_981_im; // @[Reg.scala 15:16]
  reg [31:0] out1D1_re; // @[FFT.scala 84:23]
  reg [31:0] out1D1_im; // @[FFT.scala 84:23]
  reg [31:0] _T_988_re; // @[FFT.scala 90:22]
  reg [31:0] _T_988_im; // @[FFT.scala 90:22]
  reg [31:0] _T_989_re; // @[FFT.scala 91:22]
  reg [31:0] _T_989_im; // @[FFT.scala 91:22]
  reg [9:0] _T_990; // @[FFT.scala 92:27]
  Butterfly Butterfly ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 116:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 137:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 37:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 51:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign io_dOut1_re = _T_988_re; // @[FFT.scala 90:12]
  assign io_dOut1_im = _T_988_im; // @[FFT.scala 90:12]
  assign io_dOut2_re = _T_989_re; // @[FFT.scala 91:12]
  assign io_dOut2_im = _T_989_im; // @[FFT.scala 91:12]
  assign io_dout_valid = _T_990 == 10'h1ff; // @[FFT.scala 92:17]
  assign io_busy = cnt != 10'h0; // @[FFT.scala 68:11]
  assign Butterfly_io_in1_re = _T_408_re; // @[Butterfly.scala 117:17]
  assign Butterfly_io_in1_im = 32'sh0; // @[Butterfly.scala 117:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 118:17]
  assign Butterfly_io_in2_im = 32'sh0; // @[Butterfly.scala 118:17]
  assign Butterfly_io_wn_re = 8'hff == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_255); // @[Butterfly.scala 119:16]
  assign Butterfly_io_wn_im = 8'hff == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_1023); // @[Butterfly.scala 119:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_io_in2_re = _T_537_re; // @[Butterfly.scala 139:17]
  assign Switch_io_in2_im = _T_537_im; // @[Butterfly.scala 139:17]
  assign Switch_io_sel = cnt[7]; // @[Butterfly.scala 140:17]
  assign Butterfly_1_io_in1_re = _T_673_re; // @[Butterfly.scala 117:17]
  assign Butterfly_1_io_in1_im = _T_673_im; // @[Butterfly.scala 117:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_1_io_wn_re = 7'h7f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_1919); // @[Butterfly.scala 119:16]
  assign Butterfly_1_io_wn_im = 7'h7f == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_2303); // @[Butterfly.scala 119:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_1_io_in2_re = _T_738_re; // @[Butterfly.scala 139:17]
  assign Switch_1_io_in2_im = _T_738_im; // @[Butterfly.scala 139:17]
  assign Switch_1_io_sel = cnt[6]; // @[Butterfly.scala 140:17]
  assign Butterfly_2_io_in1_re = _T_810_re; // @[Butterfly.scala 117:17]
  assign Butterfly_2_io_in1_im = _T_810_im; // @[Butterfly.scala 117:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_2_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2751); // @[Butterfly.scala 119:16]
  assign Butterfly_2_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_2943); // @[Butterfly.scala 119:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_2_io_in2_re = _T_843_re; // @[Butterfly.scala 139:17]
  assign Switch_2_io_in2_im = _T_843_im; // @[Butterfly.scala 139:17]
  assign Switch_2_io_sel = cnt[5]; // @[Butterfly.scala 140:17]
  assign Butterfly_3_io_in1_re = _T_883_re; // @[Butterfly.scala 117:17]
  assign Butterfly_3_io_in1_im = _T_883_im; // @[Butterfly.scala 117:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_3_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_3167); // @[Butterfly.scala 119:16]
  assign Butterfly_3_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_3263); // @[Butterfly.scala 119:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_3_io_in2_re = _T_900_re; // @[Butterfly.scala 139:17]
  assign Switch_3_io_in2_im = _T_900_im; // @[Butterfly.scala 139:17]
  assign Switch_3_io_sel = cnt[4]; // @[Butterfly.scala 140:17]
  assign Butterfly_4_io_in1_re = _T_924_re; // @[Butterfly.scala 117:17]
  assign Butterfly_4_io_in1_im = _T_924_im; // @[Butterfly.scala 117:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_4_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_3375); // @[Butterfly.scala 119:16]
  assign Butterfly_4_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_3423); // @[Butterfly.scala 119:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_4_io_in2_re = _T_933_re; // @[Butterfly.scala 139:17]
  assign Switch_4_io_in2_im = _T_933_im; // @[Butterfly.scala 139:17]
  assign Switch_4_io_sel = cnt[3]; // @[Butterfly.scala 140:17]
  assign Butterfly_5_io_in1_re = _T_949_re; // @[Butterfly.scala 117:17]
  assign Butterfly_5_io_in1_im = _T_949_im; // @[Butterfly.scala 117:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_5_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_3479); // @[Butterfly.scala 119:16]
  assign Butterfly_5_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_3503); // @[Butterfly.scala 119:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_5_io_in2_re = _T_954_re; // @[Butterfly.scala 139:17]
  assign Switch_5_io_in2_im = _T_954_im; // @[Butterfly.scala 139:17]
  assign Switch_5_io_sel = cnt[2]; // @[Butterfly.scala 140:17]
  assign Butterfly_6_io_in1_re = _T_966_re; // @[Butterfly.scala 117:17]
  assign Butterfly_6_io_in1_im = _T_966_im; // @[Butterfly.scala 117:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_6_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_3531); // @[Butterfly.scala 119:16]
  assign Butterfly_6_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_3543); // @[Butterfly.scala 119:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_6_io_in2_re = _T_969_re; // @[Butterfly.scala 139:17]
  assign Switch_6_io_in2_im = _T_969_im; // @[Butterfly.scala 139:17]
  assign Switch_6_io_sel = cnt[1]; // @[Butterfly.scala 140:17]
  assign Butterfly_7_io_in1_re = _T_979_re; // @[Butterfly.scala 117:17]
  assign Butterfly_7_io_in1_im = _T_979_im; // @[Butterfly.scala 117:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 118:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 118:17]
  assign Butterfly_7_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 119:16]
  assign Butterfly_7_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 119:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 138:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 138:17]
  assign Switch_7_io_in2_re = _T_981_re; // @[Butterfly.scala 139:17]
  assign Switch_7_io_in2_im = _T_981_im; // @[Butterfly.scala 139:17]
  assign Switch_7_io_sel = cnt[0]; // @[Butterfly.scala 140:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 38:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 38:17]
  assign ComplexAdd_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 39:17]
  assign ComplexAdd_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 39:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 52:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 52:17]
  assign ComplexSub_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 53:17]
  assign ComplexSub_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 53:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_153_re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_154_re = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_155_re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _T_156_re = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  _T_157_re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_158_re = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _T_159_re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_160_re = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _T_161_re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _T_162_re = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _T_163_re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _T_164_re = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  _T_165_re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _T_166_re = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  _T_167_re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  _T_168_re = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  _T_169_re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  _T_170_re = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  _T_171_re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  _T_172_re = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  _T_173_re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  _T_174_re = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  _T_175_re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  _T_176_re = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  _T_177_re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  _T_178_re = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  _T_179_re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  _T_180_re = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  _T_181_re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  _T_182_re = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  _T_183_re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  _T_184_re = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  _T_185_re = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  _T_186_re = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  _T_187_re = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  _T_188_re = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  _T_189_re = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  _T_190_re = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  _T_191_re = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  _T_192_re = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  _T_193_re = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  _T_194_re = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  _T_195_re = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  _T_196_re = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  _T_197_re = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  _T_198_re = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  _T_199_re = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  _T_200_re = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  _T_201_re = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  _T_202_re = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  _T_203_re = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  _T_204_re = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  _T_205_re = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  _T_206_re = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  _T_207_re = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  _T_208_re = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  _T_209_re = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  _T_210_re = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  _T_211_re = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  _T_212_re = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  _T_213_re = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  _T_214_re = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  _T_215_re = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  _T_216_re = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  _T_217_re = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  _T_218_re = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  _T_219_re = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  _T_220_re = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  _T_221_re = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  _T_222_re = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  _T_223_re = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  _T_224_re = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  _T_225_re = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  _T_226_re = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  _T_227_re = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  _T_228_re = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  _T_229_re = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  _T_230_re = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  _T_231_re = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  _T_232_re = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  _T_233_re = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  _T_234_re = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  _T_235_re = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  _T_236_re = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  _T_237_re = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  _T_238_re = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  _T_239_re = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  _T_240_re = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  _T_241_re = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  _T_242_re = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  _T_243_re = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  _T_244_re = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  _T_245_re = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  _T_246_re = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  _T_247_re = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  _T_248_re = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  _T_249_re = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  _T_250_re = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  _T_251_re = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  _T_252_re = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  _T_253_re = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  _T_254_re = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  _T_255_re = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  _T_256_re = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  _T_257_re = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  _T_258_re = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  _T_259_re = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  _T_260_re = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  _T_261_re = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  _T_262_re = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  _T_263_re = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  _T_264_re = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  _T_265_re = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  _T_266_re = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  _T_267_re = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  _T_268_re = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  _T_269_re = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  _T_270_re = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  _T_271_re = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  _T_272_re = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  _T_273_re = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  _T_274_re = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  _T_275_re = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  _T_276_re = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  _T_277_re = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  _T_278_re = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  _T_279_re = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  _T_280_re = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  _T_281_re = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  _T_282_re = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  _T_283_re = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  _T_284_re = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  _T_285_re = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  _T_286_re = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  _T_287_re = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  _T_288_re = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  _T_289_re = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  _T_290_re = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  _T_291_re = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  _T_292_re = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  _T_293_re = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  _T_294_re = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  _T_295_re = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  _T_296_re = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  _T_297_re = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  _T_298_re = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  _T_299_re = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  _T_300_re = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  _T_301_re = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  _T_302_re = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  _T_303_re = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  _T_304_re = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  _T_305_re = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  _T_306_re = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  _T_307_re = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  _T_308_re = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  _T_309_re = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  _T_310_re = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  _T_311_re = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  _T_312_re = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  _T_313_re = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  _T_314_re = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  _T_315_re = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  _T_316_re = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  _T_317_re = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  _T_318_re = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  _T_319_re = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  _T_320_re = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  _T_321_re = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  _T_322_re = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  _T_323_re = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  _T_324_re = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  _T_325_re = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  _T_326_re = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  _T_327_re = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  _T_328_re = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  _T_329_re = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  _T_330_re = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  _T_331_re = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  _T_332_re = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  _T_333_re = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  _T_334_re = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  _T_335_re = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  _T_336_re = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  _T_337_re = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  _T_338_re = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  _T_339_re = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  _T_340_re = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  _T_341_re = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  _T_342_re = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  _T_343_re = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  _T_344_re = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  _T_345_re = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  _T_346_re = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  _T_347_re = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  _T_348_re = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  _T_349_re = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  _T_350_re = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  _T_351_re = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  _T_352_re = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  _T_353_re = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  _T_354_re = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  _T_355_re = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  _T_356_re = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  _T_357_re = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  _T_358_re = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  _T_359_re = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  _T_360_re = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  _T_361_re = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  _T_362_re = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  _T_363_re = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  _T_364_re = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  _T_365_re = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  _T_366_re = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  _T_367_re = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  _T_368_re = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  _T_369_re = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  _T_370_re = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  _T_371_re = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  _T_372_re = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  _T_373_re = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  _T_374_re = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  _T_375_re = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  _T_376_re = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  _T_377_re = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  _T_378_re = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  _T_379_re = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  _T_380_re = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  _T_381_re = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  _T_382_re = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  _T_383_re = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  _T_384_re = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  _T_385_re = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  _T_386_re = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  _T_387_re = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  _T_388_re = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  _T_389_re = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  _T_390_re = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  _T_391_re = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  _T_392_re = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  _T_393_re = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  _T_394_re = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  _T_395_re = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  _T_396_re = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  _T_397_re = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  _T_398_re = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  _T_399_re = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  _T_400_re = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  _T_401_re = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  _T_402_re = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  _T_403_re = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  _T_404_re = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  _T_405_re = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  _T_406_re = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  _T_407_re = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  _T_408_re = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  _T_410_re = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  _T_410_im = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  _T_411_re = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  _T_411_im = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  _T_412_re = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  _T_412_im = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  _T_413_re = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  _T_413_im = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  _T_414_re = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  _T_414_im = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  _T_415_re = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  _T_415_im = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  _T_416_re = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  _T_416_im = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  _T_417_re = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  _T_417_im = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  _T_418_re = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  _T_418_im = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  _T_419_re = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  _T_419_im = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  _T_420_re = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  _T_420_im = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  _T_421_re = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  _T_421_im = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  _T_422_re = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  _T_422_im = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  _T_423_re = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  _T_423_im = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  _T_424_re = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  _T_424_im = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  _T_425_re = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  _T_425_im = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  _T_426_re = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  _T_426_im = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  _T_427_re = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  _T_427_im = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  _T_428_re = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  _T_428_im = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  _T_429_re = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  _T_429_im = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  _T_430_re = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  _T_430_im = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  _T_431_re = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  _T_431_im = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  _T_432_re = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  _T_432_im = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  _T_433_re = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  _T_433_im = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  _T_434_re = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  _T_434_im = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  _T_435_re = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  _T_435_im = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  _T_436_re = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  _T_436_im = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  _T_437_re = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  _T_437_im = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  _T_438_re = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  _T_438_im = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  _T_439_re = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  _T_439_im = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  _T_440_re = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  _T_440_im = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  _T_441_re = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  _T_441_im = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  _T_442_re = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  _T_442_im = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  _T_443_re = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  _T_443_im = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  _T_444_re = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  _T_444_im = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  _T_445_re = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  _T_445_im = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  _T_446_re = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  _T_446_im = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  _T_447_re = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  _T_447_im = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  _T_448_re = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  _T_448_im = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  _T_449_re = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  _T_449_im = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  _T_450_re = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  _T_450_im = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  _T_451_re = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  _T_451_im = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  _T_452_re = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  _T_452_im = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  _T_453_re = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  _T_453_im = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  _T_454_re = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  _T_454_im = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  _T_455_re = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  _T_455_im = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  _T_456_re = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  _T_456_im = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  _T_457_re = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  _T_457_im = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  _T_458_re = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  _T_458_im = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  _T_459_re = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  _T_459_im = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  _T_460_re = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  _T_460_im = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  _T_461_re = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  _T_461_im = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  _T_462_re = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  _T_462_im = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  _T_463_re = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  _T_463_im = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  _T_464_re = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  _T_464_im = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  _T_465_re = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  _T_465_im = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  _T_466_re = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  _T_466_im = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  _T_467_re = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  _T_467_im = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  _T_468_re = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  _T_468_im = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  _T_469_re = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  _T_469_im = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  _T_470_re = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  _T_470_im = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  _T_471_re = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  _T_471_im = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  _T_472_re = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  _T_472_im = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  _T_473_re = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  _T_473_im = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  _T_474_re = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  _T_474_im = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  _T_475_re = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  _T_475_im = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  _T_476_re = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  _T_476_im = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  _T_477_re = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  _T_477_im = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  _T_478_re = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  _T_478_im = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  _T_479_re = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  _T_479_im = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  _T_480_re = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  _T_480_im = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  _T_481_re = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  _T_481_im = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  _T_482_re = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  _T_482_im = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  _T_483_re = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  _T_483_im = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  _T_484_re = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  _T_484_im = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  _T_485_re = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  _T_485_im = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  _T_486_re = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  _T_486_im = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  _T_487_re = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  _T_487_im = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  _T_488_re = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  _T_488_im = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  _T_489_re = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  _T_489_im = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  _T_490_re = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  _T_490_im = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  _T_491_re = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  _T_491_im = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  _T_492_re = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  _T_492_im = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  _T_493_re = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  _T_493_im = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  _T_494_re = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  _T_494_im = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  _T_495_re = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  _T_495_im = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  _T_496_re = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  _T_496_im = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  _T_497_re = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  _T_497_im = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  _T_498_re = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  _T_498_im = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  _T_499_re = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  _T_499_im = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  _T_500_re = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  _T_500_im = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  _T_501_re = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  _T_501_im = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  _T_502_re = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  _T_502_im = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  _T_503_re = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  _T_503_im = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  _T_504_re = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  _T_504_im = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  _T_505_re = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  _T_505_im = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  _T_506_re = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  _T_506_im = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  _T_507_re = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  _T_507_im = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  _T_508_re = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  _T_508_im = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  _T_509_re = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  _T_509_im = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  _T_510_re = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  _T_510_im = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  _T_511_re = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  _T_511_im = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  _T_512_re = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  _T_512_im = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  _T_513_re = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  _T_513_im = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  _T_514_re = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  _T_514_im = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  _T_515_re = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  _T_515_im = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  _T_516_re = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  _T_516_im = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  _T_517_re = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  _T_517_im = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  _T_518_re = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  _T_518_im = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  _T_519_re = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  _T_519_im = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  _T_520_re = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  _T_520_im = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  _T_521_re = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  _T_521_im = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  _T_522_re = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  _T_522_im = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  _T_523_re = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  _T_523_im = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  _T_524_re = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  _T_524_im = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  _T_525_re = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  _T_525_im = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  _T_526_re = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  _T_526_im = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  _T_527_re = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  _T_527_im = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  _T_528_re = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  _T_528_im = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  _T_529_re = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  _T_529_im = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  _T_530_re = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  _T_530_im = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  _T_531_re = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  _T_531_im = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  _T_532_re = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  _T_532_im = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  _T_533_re = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  _T_533_im = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  _T_534_re = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  _T_534_im = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  _T_535_re = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  _T_535_im = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  _T_536_re = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  _T_536_im = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  _T_537_re = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  _T_537_im = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  _T_546_re = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  _T_546_im = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  _T_547_re = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  _T_547_im = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  _T_548_re = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  _T_548_im = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  _T_549_re = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  _T_549_im = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  _T_550_re = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  _T_550_im = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  _T_551_re = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  _T_551_im = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  _T_552_re = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  _T_552_im = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  _T_553_re = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  _T_553_im = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  _T_554_re = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  _T_554_im = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  _T_555_re = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  _T_555_im = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  _T_556_re = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  _T_556_im = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  _T_557_re = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  _T_557_im = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  _T_558_re = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  _T_558_im = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  _T_559_re = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  _T_559_im = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  _T_560_re = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  _T_560_im = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  _T_561_re = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  _T_561_im = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  _T_562_re = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  _T_562_im = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  _T_563_re = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  _T_563_im = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  _T_564_re = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  _T_564_im = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  _T_565_re = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  _T_565_im = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  _T_566_re = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  _T_566_im = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  _T_567_re = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  _T_567_im = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  _T_568_re = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  _T_568_im = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  _T_569_re = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  _T_569_im = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  _T_570_re = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  _T_570_im = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  _T_571_re = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  _T_571_im = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  _T_572_re = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  _T_572_im = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  _T_573_re = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  _T_573_im = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  _T_574_re = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  _T_574_im = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  _T_575_re = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  _T_575_im = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  _T_576_re = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  _T_576_im = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  _T_577_re = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  _T_577_im = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  _T_578_re = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  _T_578_im = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  _T_579_re = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  _T_579_im = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  _T_580_re = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  _T_580_im = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  _T_581_re = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  _T_581_im = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  _T_582_re = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  _T_582_im = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  _T_583_re = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  _T_583_im = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  _T_584_re = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  _T_584_im = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  _T_585_re = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  _T_585_im = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  _T_586_re = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  _T_586_im = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  _T_587_re = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  _T_587_im = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  _T_588_re = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  _T_588_im = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  _T_589_re = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  _T_589_im = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  _T_590_re = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  _T_590_im = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  _T_591_re = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  _T_591_im = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  _T_592_re = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  _T_592_im = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  _T_593_re = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  _T_593_im = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  _T_594_re = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  _T_594_im = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  _T_595_re = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  _T_595_im = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  _T_596_re = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  _T_596_im = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  _T_597_re = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  _T_597_im = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  _T_598_re = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  _T_598_im = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  _T_599_re = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  _T_599_im = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  _T_600_re = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  _T_600_im = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  _T_601_re = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  _T_601_im = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  _T_602_re = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  _T_602_im = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  _T_603_re = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  _T_603_im = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  _T_604_re = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  _T_604_im = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  _T_605_re = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  _T_605_im = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  _T_606_re = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  _T_606_im = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  _T_607_re = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  _T_607_im = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  _T_608_re = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  _T_608_im = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  _T_609_re = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  _T_609_im = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  _T_610_re = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  _T_610_im = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  _T_611_re = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  _T_611_im = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  _T_612_re = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  _T_612_im = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  _T_613_re = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  _T_613_im = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  _T_614_re = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  _T_614_im = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  _T_615_re = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  _T_615_im = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  _T_616_re = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  _T_616_im = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  _T_617_re = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  _T_617_im = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  _T_618_re = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  _T_618_im = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  _T_619_re = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  _T_619_im = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  _T_620_re = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  _T_620_im = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  _T_621_re = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  _T_621_im = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  _T_622_re = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  _T_622_im = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  _T_623_re = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  _T_623_im = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  _T_624_re = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  _T_624_im = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  _T_625_re = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  _T_625_im = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  _T_626_re = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  _T_626_im = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  _T_627_re = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  _T_627_im = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  _T_628_re = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  _T_628_im = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  _T_629_re = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  _T_629_im = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  _T_630_re = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  _T_630_im = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  _T_631_re = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  _T_631_im = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  _T_632_re = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  _T_632_im = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  _T_633_re = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  _T_633_im = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  _T_634_re = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  _T_634_im = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  _T_635_re = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  _T_635_im = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  _T_636_re = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  _T_636_im = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  _T_637_re = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  _T_637_im = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  _T_638_re = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  _T_638_im = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  _T_639_re = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  _T_639_im = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  _T_640_re = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  _T_640_im = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  _T_641_re = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  _T_641_im = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  _T_642_re = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  _T_642_im = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  _T_643_re = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  _T_643_im = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  _T_644_re = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  _T_644_im = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  _T_645_re = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  _T_645_im = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  _T_646_re = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  _T_646_im = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  _T_647_re = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  _T_647_im = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  _T_648_re = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  _T_648_im = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  _T_649_re = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  _T_649_im = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  _T_650_re = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  _T_650_im = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  _T_651_re = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  _T_651_im = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  _T_652_re = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  _T_652_im = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  _T_653_re = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  _T_653_im = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  _T_654_re = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  _T_654_im = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  _T_655_re = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  _T_655_im = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  _T_656_re = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  _T_656_im = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  _T_657_re = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  _T_657_im = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  _T_658_re = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  _T_658_im = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  _T_659_re = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  _T_659_im = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  _T_660_re = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  _T_660_im = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  _T_661_re = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  _T_661_im = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  _T_662_re = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  _T_662_im = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  _T_663_re = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  _T_663_im = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  _T_664_re = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  _T_664_im = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  _T_665_re = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  _T_665_im = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  _T_666_re = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  _T_666_im = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  _T_667_re = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  _T_667_im = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  _T_668_re = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  _T_668_im = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  _T_669_re = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  _T_669_im = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  _T_670_re = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  _T_670_im = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  _T_671_re = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  _T_671_im = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  _T_672_re = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  _T_672_im = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  _T_673_re = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  _T_673_im = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  _T_675_re = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  _T_675_im = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  _T_676_re = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  _T_676_im = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  _T_677_re = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  _T_677_im = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  _T_678_re = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  _T_678_im = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  _T_679_re = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  _T_679_im = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  _T_680_re = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  _T_680_im = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  _T_681_re = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  _T_681_im = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  _T_682_re = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  _T_682_im = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  _T_683_re = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  _T_683_im = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  _T_684_re = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  _T_684_im = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  _T_685_re = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  _T_685_im = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  _T_686_re = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  _T_686_im = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  _T_687_re = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  _T_687_im = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  _T_688_re = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  _T_688_im = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  _T_689_re = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  _T_689_im = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  _T_690_re = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  _T_690_im = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  _T_691_re = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  _T_691_im = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  _T_692_re = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  _T_692_im = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  _T_693_re = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  _T_693_im = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  _T_694_re = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  _T_694_im = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  _T_695_re = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  _T_695_im = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  _T_696_re = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  _T_696_im = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  _T_697_re = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  _T_697_im = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  _T_698_re = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  _T_698_im = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  _T_699_re = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  _T_699_im = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  _T_700_re = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  _T_700_im = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  _T_701_re = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  _T_701_im = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  _T_702_re = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  _T_702_im = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  _T_703_re = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  _T_703_im = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  _T_704_re = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  _T_704_im = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  _T_705_re = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  _T_705_im = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  _T_706_re = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  _T_706_im = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  _T_707_re = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  _T_707_im = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  _T_708_re = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  _T_708_im = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  _T_709_re = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  _T_709_im = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  _T_710_re = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  _T_710_im = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  _T_711_re = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  _T_711_im = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  _T_712_re = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  _T_712_im = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  _T_713_re = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  _T_713_im = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  _T_714_re = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  _T_714_im = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  _T_715_re = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  _T_715_im = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  _T_716_re = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  _T_716_im = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  _T_717_re = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  _T_717_im = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  _T_718_re = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  _T_718_im = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  _T_719_re = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  _T_719_im = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  _T_720_re = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  _T_720_im = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  _T_721_re = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  _T_721_im = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  _T_722_re = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  _T_722_im = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  _T_723_re = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  _T_723_im = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  _T_724_re = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  _T_724_im = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  _T_725_re = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  _T_725_im = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  _T_726_re = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  _T_726_im = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  _T_727_re = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  _T_727_im = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  _T_728_re = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  _T_728_im = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  _T_729_re = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  _T_729_im = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  _T_730_re = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  _T_730_im = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  _T_731_re = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  _T_731_im = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  _T_732_re = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  _T_732_im = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  _T_733_re = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  _T_733_im = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  _T_734_re = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  _T_734_im = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  _T_735_re = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  _T_735_im = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  _T_736_re = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  _T_736_im = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  _T_737_re = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  _T_737_im = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  _T_738_re = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  _T_738_im = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  _T_747_re = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  _T_747_im = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  _T_748_re = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  _T_748_im = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  _T_749_re = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  _T_749_im = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  _T_750_re = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  _T_750_im = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  _T_751_re = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  _T_751_im = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  _T_752_re = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  _T_752_im = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  _T_753_re = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  _T_753_im = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  _T_754_re = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  _T_754_im = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  _T_755_re = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  _T_755_im = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  _T_756_re = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  _T_756_im = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  _T_757_re = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  _T_757_im = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  _T_758_re = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  _T_758_im = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  _T_759_re = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  _T_759_im = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  _T_760_re = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  _T_760_im = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  _T_761_re = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  _T_761_im = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  _T_762_re = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  _T_762_im = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  _T_763_re = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  _T_763_im = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  _T_764_re = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  _T_764_im = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  _T_765_re = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  _T_765_im = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  _T_766_re = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  _T_766_im = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  _T_767_re = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  _T_767_im = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  _T_768_re = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  _T_768_im = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  _T_769_re = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  _T_769_im = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  _T_770_re = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  _T_770_im = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  _T_771_re = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  _T_771_im = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  _T_772_re = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  _T_772_im = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  _T_773_re = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  _T_773_im = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  _T_774_re = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  _T_774_im = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  _T_775_re = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  _T_775_im = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  _T_776_re = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  _T_776_im = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  _T_777_re = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  _T_777_im = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  _T_778_re = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  _T_778_im = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  _T_779_re = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  _T_779_im = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  _T_780_re = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  _T_780_im = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  _T_781_re = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  _T_781_im = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  _T_782_re = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  _T_782_im = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  _T_783_re = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  _T_783_im = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  _T_784_re = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  _T_784_im = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  _T_785_re = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  _T_785_im = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  _T_786_re = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  _T_786_im = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  _T_787_re = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  _T_787_im = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  _T_788_re = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  _T_788_im = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  _T_789_re = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  _T_789_im = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  _T_790_re = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  _T_790_im = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  _T_791_re = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  _T_791_im = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  _T_792_re = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  _T_792_im = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  _T_793_re = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  _T_793_im = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  _T_794_re = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  _T_794_im = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  _T_795_re = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  _T_795_im = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  _T_796_re = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  _T_796_im = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  _T_797_re = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  _T_797_im = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  _T_798_re = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  _T_798_im = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  _T_799_re = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  _T_799_im = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  _T_800_re = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  _T_800_im = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  _T_801_re = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  _T_801_im = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  _T_802_re = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  _T_802_im = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  _T_803_re = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  _T_803_im = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  _T_804_re = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  _T_804_im = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  _T_805_re = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  _T_805_im = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  _T_806_re = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  _T_806_im = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  _T_807_re = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  _T_807_im = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  _T_808_re = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  _T_808_im = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  _T_809_re = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  _T_809_im = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  _T_810_re = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  _T_810_im = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  _T_812_re = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  _T_812_im = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  _T_813_re = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  _T_813_im = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  _T_814_re = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  _T_814_im = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  _T_815_re = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  _T_815_im = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  _T_816_re = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  _T_816_im = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  _T_817_re = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  _T_817_im = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  _T_818_re = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  _T_818_im = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  _T_819_re = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  _T_819_im = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  _T_820_re = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  _T_820_im = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  _T_821_re = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  _T_821_im = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  _T_822_re = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  _T_822_im = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  _T_823_re = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  _T_823_im = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  _T_824_re = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  _T_824_im = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  _T_825_re = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  _T_825_im = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  _T_826_re = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  _T_826_im = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  _T_827_re = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  _T_827_im = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  _T_828_re = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  _T_828_im = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  _T_829_re = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  _T_829_im = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  _T_830_re = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  _T_830_im = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  _T_831_re = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  _T_831_im = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  _T_832_re = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  _T_832_im = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  _T_833_re = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  _T_833_im = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  _T_834_re = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  _T_834_im = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  _T_835_re = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  _T_835_im = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  _T_836_re = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  _T_836_im = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  _T_837_re = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  _T_837_im = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  _T_838_re = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  _T_838_im = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  _T_839_re = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  _T_839_im = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  _T_840_re = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  _T_840_im = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  _T_841_re = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  _T_841_im = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  _T_842_re = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  _T_842_im = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  _T_843_re = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  _T_843_im = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  _T_852_re = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  _T_852_im = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  _T_853_re = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  _T_853_im = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  _T_854_re = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  _T_854_im = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  _T_855_re = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  _T_855_im = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  _T_856_re = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  _T_856_im = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  _T_857_re = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  _T_857_im = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  _T_858_re = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  _T_858_im = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  _T_859_re = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  _T_859_im = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  _T_860_re = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  _T_860_im = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  _T_861_re = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  _T_861_im = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  _T_862_re = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  _T_862_im = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  _T_863_re = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  _T_863_im = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  _T_864_re = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  _T_864_im = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  _T_865_re = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  _T_865_im = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  _T_866_re = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  _T_866_im = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  _T_867_re = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  _T_867_im = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  _T_868_re = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  _T_868_im = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  _T_869_re = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  _T_869_im = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  _T_870_re = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  _T_870_im = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  _T_871_re = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  _T_871_im = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  _T_872_re = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  _T_872_im = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  _T_873_re = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  _T_873_im = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  _T_874_re = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  _T_874_im = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  _T_875_re = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  _T_875_im = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  _T_876_re = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  _T_876_im = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  _T_877_re = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  _T_877_im = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  _T_878_re = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  _T_878_im = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  _T_879_re = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  _T_879_im = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  _T_880_re = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  _T_880_im = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  _T_881_re = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  _T_881_im = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  _T_882_re = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  _T_882_im = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  _T_883_re = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  _T_883_im = _RAND_1152[31:0];
  _RAND_1153 = {1{`RANDOM}};
  _T_885_re = _RAND_1153[31:0];
  _RAND_1154 = {1{`RANDOM}};
  _T_885_im = _RAND_1154[31:0];
  _RAND_1155 = {1{`RANDOM}};
  _T_886_re = _RAND_1155[31:0];
  _RAND_1156 = {1{`RANDOM}};
  _T_886_im = _RAND_1156[31:0];
  _RAND_1157 = {1{`RANDOM}};
  _T_887_re = _RAND_1157[31:0];
  _RAND_1158 = {1{`RANDOM}};
  _T_887_im = _RAND_1158[31:0];
  _RAND_1159 = {1{`RANDOM}};
  _T_888_re = _RAND_1159[31:0];
  _RAND_1160 = {1{`RANDOM}};
  _T_888_im = _RAND_1160[31:0];
  _RAND_1161 = {1{`RANDOM}};
  _T_889_re = _RAND_1161[31:0];
  _RAND_1162 = {1{`RANDOM}};
  _T_889_im = _RAND_1162[31:0];
  _RAND_1163 = {1{`RANDOM}};
  _T_890_re = _RAND_1163[31:0];
  _RAND_1164 = {1{`RANDOM}};
  _T_890_im = _RAND_1164[31:0];
  _RAND_1165 = {1{`RANDOM}};
  _T_891_re = _RAND_1165[31:0];
  _RAND_1166 = {1{`RANDOM}};
  _T_891_im = _RAND_1166[31:0];
  _RAND_1167 = {1{`RANDOM}};
  _T_892_re = _RAND_1167[31:0];
  _RAND_1168 = {1{`RANDOM}};
  _T_892_im = _RAND_1168[31:0];
  _RAND_1169 = {1{`RANDOM}};
  _T_893_re = _RAND_1169[31:0];
  _RAND_1170 = {1{`RANDOM}};
  _T_893_im = _RAND_1170[31:0];
  _RAND_1171 = {1{`RANDOM}};
  _T_894_re = _RAND_1171[31:0];
  _RAND_1172 = {1{`RANDOM}};
  _T_894_im = _RAND_1172[31:0];
  _RAND_1173 = {1{`RANDOM}};
  _T_895_re = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  _T_895_im = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  _T_896_re = _RAND_1175[31:0];
  _RAND_1176 = {1{`RANDOM}};
  _T_896_im = _RAND_1176[31:0];
  _RAND_1177 = {1{`RANDOM}};
  _T_897_re = _RAND_1177[31:0];
  _RAND_1178 = {1{`RANDOM}};
  _T_897_im = _RAND_1178[31:0];
  _RAND_1179 = {1{`RANDOM}};
  _T_898_re = _RAND_1179[31:0];
  _RAND_1180 = {1{`RANDOM}};
  _T_898_im = _RAND_1180[31:0];
  _RAND_1181 = {1{`RANDOM}};
  _T_899_re = _RAND_1181[31:0];
  _RAND_1182 = {1{`RANDOM}};
  _T_899_im = _RAND_1182[31:0];
  _RAND_1183 = {1{`RANDOM}};
  _T_900_re = _RAND_1183[31:0];
  _RAND_1184 = {1{`RANDOM}};
  _T_900_im = _RAND_1184[31:0];
  _RAND_1185 = {1{`RANDOM}};
  _T_909_re = _RAND_1185[31:0];
  _RAND_1186 = {1{`RANDOM}};
  _T_909_im = _RAND_1186[31:0];
  _RAND_1187 = {1{`RANDOM}};
  _T_910_re = _RAND_1187[31:0];
  _RAND_1188 = {1{`RANDOM}};
  _T_910_im = _RAND_1188[31:0];
  _RAND_1189 = {1{`RANDOM}};
  _T_911_re = _RAND_1189[31:0];
  _RAND_1190 = {1{`RANDOM}};
  _T_911_im = _RAND_1190[31:0];
  _RAND_1191 = {1{`RANDOM}};
  _T_912_re = _RAND_1191[31:0];
  _RAND_1192 = {1{`RANDOM}};
  _T_912_im = _RAND_1192[31:0];
  _RAND_1193 = {1{`RANDOM}};
  _T_913_re = _RAND_1193[31:0];
  _RAND_1194 = {1{`RANDOM}};
  _T_913_im = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  _T_914_re = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  _T_914_im = _RAND_1196[31:0];
  _RAND_1197 = {1{`RANDOM}};
  _T_915_re = _RAND_1197[31:0];
  _RAND_1198 = {1{`RANDOM}};
  _T_915_im = _RAND_1198[31:0];
  _RAND_1199 = {1{`RANDOM}};
  _T_916_re = _RAND_1199[31:0];
  _RAND_1200 = {1{`RANDOM}};
  _T_916_im = _RAND_1200[31:0];
  _RAND_1201 = {1{`RANDOM}};
  _T_917_re = _RAND_1201[31:0];
  _RAND_1202 = {1{`RANDOM}};
  _T_917_im = _RAND_1202[31:0];
  _RAND_1203 = {1{`RANDOM}};
  _T_918_re = _RAND_1203[31:0];
  _RAND_1204 = {1{`RANDOM}};
  _T_918_im = _RAND_1204[31:0];
  _RAND_1205 = {1{`RANDOM}};
  _T_919_re = _RAND_1205[31:0];
  _RAND_1206 = {1{`RANDOM}};
  _T_919_im = _RAND_1206[31:0];
  _RAND_1207 = {1{`RANDOM}};
  _T_920_re = _RAND_1207[31:0];
  _RAND_1208 = {1{`RANDOM}};
  _T_920_im = _RAND_1208[31:0];
  _RAND_1209 = {1{`RANDOM}};
  _T_921_re = _RAND_1209[31:0];
  _RAND_1210 = {1{`RANDOM}};
  _T_921_im = _RAND_1210[31:0];
  _RAND_1211 = {1{`RANDOM}};
  _T_922_re = _RAND_1211[31:0];
  _RAND_1212 = {1{`RANDOM}};
  _T_922_im = _RAND_1212[31:0];
  _RAND_1213 = {1{`RANDOM}};
  _T_923_re = _RAND_1213[31:0];
  _RAND_1214 = {1{`RANDOM}};
  _T_923_im = _RAND_1214[31:0];
  _RAND_1215 = {1{`RANDOM}};
  _T_924_re = _RAND_1215[31:0];
  _RAND_1216 = {1{`RANDOM}};
  _T_924_im = _RAND_1216[31:0];
  _RAND_1217 = {1{`RANDOM}};
  _T_926_re = _RAND_1217[31:0];
  _RAND_1218 = {1{`RANDOM}};
  _T_926_im = _RAND_1218[31:0];
  _RAND_1219 = {1{`RANDOM}};
  _T_927_re = _RAND_1219[31:0];
  _RAND_1220 = {1{`RANDOM}};
  _T_927_im = _RAND_1220[31:0];
  _RAND_1221 = {1{`RANDOM}};
  _T_928_re = _RAND_1221[31:0];
  _RAND_1222 = {1{`RANDOM}};
  _T_928_im = _RAND_1222[31:0];
  _RAND_1223 = {1{`RANDOM}};
  _T_929_re = _RAND_1223[31:0];
  _RAND_1224 = {1{`RANDOM}};
  _T_929_im = _RAND_1224[31:0];
  _RAND_1225 = {1{`RANDOM}};
  _T_930_re = _RAND_1225[31:0];
  _RAND_1226 = {1{`RANDOM}};
  _T_930_im = _RAND_1226[31:0];
  _RAND_1227 = {1{`RANDOM}};
  _T_931_re = _RAND_1227[31:0];
  _RAND_1228 = {1{`RANDOM}};
  _T_931_im = _RAND_1228[31:0];
  _RAND_1229 = {1{`RANDOM}};
  _T_932_re = _RAND_1229[31:0];
  _RAND_1230 = {1{`RANDOM}};
  _T_932_im = _RAND_1230[31:0];
  _RAND_1231 = {1{`RANDOM}};
  _T_933_re = _RAND_1231[31:0];
  _RAND_1232 = {1{`RANDOM}};
  _T_933_im = _RAND_1232[31:0];
  _RAND_1233 = {1{`RANDOM}};
  _T_942_re = _RAND_1233[31:0];
  _RAND_1234 = {1{`RANDOM}};
  _T_942_im = _RAND_1234[31:0];
  _RAND_1235 = {1{`RANDOM}};
  _T_943_re = _RAND_1235[31:0];
  _RAND_1236 = {1{`RANDOM}};
  _T_943_im = _RAND_1236[31:0];
  _RAND_1237 = {1{`RANDOM}};
  _T_944_re = _RAND_1237[31:0];
  _RAND_1238 = {1{`RANDOM}};
  _T_944_im = _RAND_1238[31:0];
  _RAND_1239 = {1{`RANDOM}};
  _T_945_re = _RAND_1239[31:0];
  _RAND_1240 = {1{`RANDOM}};
  _T_945_im = _RAND_1240[31:0];
  _RAND_1241 = {1{`RANDOM}};
  _T_946_re = _RAND_1241[31:0];
  _RAND_1242 = {1{`RANDOM}};
  _T_946_im = _RAND_1242[31:0];
  _RAND_1243 = {1{`RANDOM}};
  _T_947_re = _RAND_1243[31:0];
  _RAND_1244 = {1{`RANDOM}};
  _T_947_im = _RAND_1244[31:0];
  _RAND_1245 = {1{`RANDOM}};
  _T_948_re = _RAND_1245[31:0];
  _RAND_1246 = {1{`RANDOM}};
  _T_948_im = _RAND_1246[31:0];
  _RAND_1247 = {1{`RANDOM}};
  _T_949_re = _RAND_1247[31:0];
  _RAND_1248 = {1{`RANDOM}};
  _T_949_im = _RAND_1248[31:0];
  _RAND_1249 = {1{`RANDOM}};
  _T_951_re = _RAND_1249[31:0];
  _RAND_1250 = {1{`RANDOM}};
  _T_951_im = _RAND_1250[31:0];
  _RAND_1251 = {1{`RANDOM}};
  _T_952_re = _RAND_1251[31:0];
  _RAND_1252 = {1{`RANDOM}};
  _T_952_im = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  _T_953_re = _RAND_1253[31:0];
  _RAND_1254 = {1{`RANDOM}};
  _T_953_im = _RAND_1254[31:0];
  _RAND_1255 = {1{`RANDOM}};
  _T_954_re = _RAND_1255[31:0];
  _RAND_1256 = {1{`RANDOM}};
  _T_954_im = _RAND_1256[31:0];
  _RAND_1257 = {1{`RANDOM}};
  _T_963_re = _RAND_1257[31:0];
  _RAND_1258 = {1{`RANDOM}};
  _T_963_im = _RAND_1258[31:0];
  _RAND_1259 = {1{`RANDOM}};
  _T_964_re = _RAND_1259[31:0];
  _RAND_1260 = {1{`RANDOM}};
  _T_964_im = _RAND_1260[31:0];
  _RAND_1261 = {1{`RANDOM}};
  _T_965_re = _RAND_1261[31:0];
  _RAND_1262 = {1{`RANDOM}};
  _T_965_im = _RAND_1262[31:0];
  _RAND_1263 = {1{`RANDOM}};
  _T_966_re = _RAND_1263[31:0];
  _RAND_1264 = {1{`RANDOM}};
  _T_966_im = _RAND_1264[31:0];
  _RAND_1265 = {1{`RANDOM}};
  _T_968_re = _RAND_1265[31:0];
  _RAND_1266 = {1{`RANDOM}};
  _T_968_im = _RAND_1266[31:0];
  _RAND_1267 = {1{`RANDOM}};
  _T_969_re = _RAND_1267[31:0];
  _RAND_1268 = {1{`RANDOM}};
  _T_969_im = _RAND_1268[31:0];
  _RAND_1269 = {1{`RANDOM}};
  _T_978_re = _RAND_1269[31:0];
  _RAND_1270 = {1{`RANDOM}};
  _T_978_im = _RAND_1270[31:0];
  _RAND_1271 = {1{`RANDOM}};
  _T_979_re = _RAND_1271[31:0];
  _RAND_1272 = {1{`RANDOM}};
  _T_979_im = _RAND_1272[31:0];
  _RAND_1273 = {1{`RANDOM}};
  _T_981_re = _RAND_1273[31:0];
  _RAND_1274 = {1{`RANDOM}};
  _T_981_im = _RAND_1274[31:0];
  _RAND_1275 = {1{`RANDOM}};
  out1D1_re = _RAND_1275[31:0];
  _RAND_1276 = {1{`RANDOM}};
  out1D1_im = _RAND_1276[31:0];
  _RAND_1277 = {1{`RANDOM}};
  _T_988_re = _RAND_1277[31:0];
  _RAND_1278 = {1{`RANDOM}};
  _T_988_im = _RAND_1278[31:0];
  _RAND_1279 = {1{`RANDOM}};
  _T_989_re = _RAND_1279[31:0];
  _RAND_1280 = {1{`RANDOM}};
  _T_989_im = _RAND_1280[31:0];
  _RAND_1281 = {1{`RANDOM}};
  _T_990 = _RAND_1281[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 10'h0;
    end else if (_T) begin
      if (_T_1) begin
        cnt <= 10'h0;
      end else begin
        cnt <= _T_3;
      end
    end
    _T_153_re <= io_dIn_re;
    _T_154_re <= _T_153_re;
    _T_155_re <= _T_154_re;
    _T_156_re <= _T_155_re;
    _T_157_re <= _T_156_re;
    _T_158_re <= _T_157_re;
    _T_159_re <= _T_158_re;
    _T_160_re <= _T_159_re;
    _T_161_re <= _T_160_re;
    _T_162_re <= _T_161_re;
    _T_163_re <= _T_162_re;
    _T_164_re <= _T_163_re;
    _T_165_re <= _T_164_re;
    _T_166_re <= _T_165_re;
    _T_167_re <= _T_166_re;
    _T_168_re <= _T_167_re;
    _T_169_re <= _T_168_re;
    _T_170_re <= _T_169_re;
    _T_171_re <= _T_170_re;
    _T_172_re <= _T_171_re;
    _T_173_re <= _T_172_re;
    _T_174_re <= _T_173_re;
    _T_175_re <= _T_174_re;
    _T_176_re <= _T_175_re;
    _T_177_re <= _T_176_re;
    _T_178_re <= _T_177_re;
    _T_179_re <= _T_178_re;
    _T_180_re <= _T_179_re;
    _T_181_re <= _T_180_re;
    _T_182_re <= _T_181_re;
    _T_183_re <= _T_182_re;
    _T_184_re <= _T_183_re;
    _T_185_re <= _T_184_re;
    _T_186_re <= _T_185_re;
    _T_187_re <= _T_186_re;
    _T_188_re <= _T_187_re;
    _T_189_re <= _T_188_re;
    _T_190_re <= _T_189_re;
    _T_191_re <= _T_190_re;
    _T_192_re <= _T_191_re;
    _T_193_re <= _T_192_re;
    _T_194_re <= _T_193_re;
    _T_195_re <= _T_194_re;
    _T_196_re <= _T_195_re;
    _T_197_re <= _T_196_re;
    _T_198_re <= _T_197_re;
    _T_199_re <= _T_198_re;
    _T_200_re <= _T_199_re;
    _T_201_re <= _T_200_re;
    _T_202_re <= _T_201_re;
    _T_203_re <= _T_202_re;
    _T_204_re <= _T_203_re;
    _T_205_re <= _T_204_re;
    _T_206_re <= _T_205_re;
    _T_207_re <= _T_206_re;
    _T_208_re <= _T_207_re;
    _T_209_re <= _T_208_re;
    _T_210_re <= _T_209_re;
    _T_211_re <= _T_210_re;
    _T_212_re <= _T_211_re;
    _T_213_re <= _T_212_re;
    _T_214_re <= _T_213_re;
    _T_215_re <= _T_214_re;
    _T_216_re <= _T_215_re;
    _T_217_re <= _T_216_re;
    _T_218_re <= _T_217_re;
    _T_219_re <= _T_218_re;
    _T_220_re <= _T_219_re;
    _T_221_re <= _T_220_re;
    _T_222_re <= _T_221_re;
    _T_223_re <= _T_222_re;
    _T_224_re <= _T_223_re;
    _T_225_re <= _T_224_re;
    _T_226_re <= _T_225_re;
    _T_227_re <= _T_226_re;
    _T_228_re <= _T_227_re;
    _T_229_re <= _T_228_re;
    _T_230_re <= _T_229_re;
    _T_231_re <= _T_230_re;
    _T_232_re <= _T_231_re;
    _T_233_re <= _T_232_re;
    _T_234_re <= _T_233_re;
    _T_235_re <= _T_234_re;
    _T_236_re <= _T_235_re;
    _T_237_re <= _T_236_re;
    _T_238_re <= _T_237_re;
    _T_239_re <= _T_238_re;
    _T_240_re <= _T_239_re;
    _T_241_re <= _T_240_re;
    _T_242_re <= _T_241_re;
    _T_243_re <= _T_242_re;
    _T_244_re <= _T_243_re;
    _T_245_re <= _T_244_re;
    _T_246_re <= _T_245_re;
    _T_247_re <= _T_246_re;
    _T_248_re <= _T_247_re;
    _T_249_re <= _T_248_re;
    _T_250_re <= _T_249_re;
    _T_251_re <= _T_250_re;
    _T_252_re <= _T_251_re;
    _T_253_re <= _T_252_re;
    _T_254_re <= _T_253_re;
    _T_255_re <= _T_254_re;
    _T_256_re <= _T_255_re;
    _T_257_re <= _T_256_re;
    _T_258_re <= _T_257_re;
    _T_259_re <= _T_258_re;
    _T_260_re <= _T_259_re;
    _T_261_re <= _T_260_re;
    _T_262_re <= _T_261_re;
    _T_263_re <= _T_262_re;
    _T_264_re <= _T_263_re;
    _T_265_re <= _T_264_re;
    _T_266_re <= _T_265_re;
    _T_267_re <= _T_266_re;
    _T_268_re <= _T_267_re;
    _T_269_re <= _T_268_re;
    _T_270_re <= _T_269_re;
    _T_271_re <= _T_270_re;
    _T_272_re <= _T_271_re;
    _T_273_re <= _T_272_re;
    _T_274_re <= _T_273_re;
    _T_275_re <= _T_274_re;
    _T_276_re <= _T_275_re;
    _T_277_re <= _T_276_re;
    _T_278_re <= _T_277_re;
    _T_279_re <= _T_278_re;
    _T_280_re <= _T_279_re;
    _T_281_re <= _T_280_re;
    _T_282_re <= _T_281_re;
    _T_283_re <= _T_282_re;
    _T_284_re <= _T_283_re;
    _T_285_re <= _T_284_re;
    _T_286_re <= _T_285_re;
    _T_287_re <= _T_286_re;
    _T_288_re <= _T_287_re;
    _T_289_re <= _T_288_re;
    _T_290_re <= _T_289_re;
    _T_291_re <= _T_290_re;
    _T_292_re <= _T_291_re;
    _T_293_re <= _T_292_re;
    _T_294_re <= _T_293_re;
    _T_295_re <= _T_294_re;
    _T_296_re <= _T_295_re;
    _T_297_re <= _T_296_re;
    _T_298_re <= _T_297_re;
    _T_299_re <= _T_298_re;
    _T_300_re <= _T_299_re;
    _T_301_re <= _T_300_re;
    _T_302_re <= _T_301_re;
    _T_303_re <= _T_302_re;
    _T_304_re <= _T_303_re;
    _T_305_re <= _T_304_re;
    _T_306_re <= _T_305_re;
    _T_307_re <= _T_306_re;
    _T_308_re <= _T_307_re;
    _T_309_re <= _T_308_re;
    _T_310_re <= _T_309_re;
    _T_311_re <= _T_310_re;
    _T_312_re <= _T_311_re;
    _T_313_re <= _T_312_re;
    _T_314_re <= _T_313_re;
    _T_315_re <= _T_314_re;
    _T_316_re <= _T_315_re;
    _T_317_re <= _T_316_re;
    _T_318_re <= _T_317_re;
    _T_319_re <= _T_318_re;
    _T_320_re <= _T_319_re;
    _T_321_re <= _T_320_re;
    _T_322_re <= _T_321_re;
    _T_323_re <= _T_322_re;
    _T_324_re <= _T_323_re;
    _T_325_re <= _T_324_re;
    _T_326_re <= _T_325_re;
    _T_327_re <= _T_326_re;
    _T_328_re <= _T_327_re;
    _T_329_re <= _T_328_re;
    _T_330_re <= _T_329_re;
    _T_331_re <= _T_330_re;
    _T_332_re <= _T_331_re;
    _T_333_re <= _T_332_re;
    _T_334_re <= _T_333_re;
    _T_335_re <= _T_334_re;
    _T_336_re <= _T_335_re;
    _T_337_re <= _T_336_re;
    _T_338_re <= _T_337_re;
    _T_339_re <= _T_338_re;
    _T_340_re <= _T_339_re;
    _T_341_re <= _T_340_re;
    _T_342_re <= _T_341_re;
    _T_343_re <= _T_342_re;
    _T_344_re <= _T_343_re;
    _T_345_re <= _T_344_re;
    _T_346_re <= _T_345_re;
    _T_347_re <= _T_346_re;
    _T_348_re <= _T_347_re;
    _T_349_re <= _T_348_re;
    _T_350_re <= _T_349_re;
    _T_351_re <= _T_350_re;
    _T_352_re <= _T_351_re;
    _T_353_re <= _T_352_re;
    _T_354_re <= _T_353_re;
    _T_355_re <= _T_354_re;
    _T_356_re <= _T_355_re;
    _T_357_re <= _T_356_re;
    _T_358_re <= _T_357_re;
    _T_359_re <= _T_358_re;
    _T_360_re <= _T_359_re;
    _T_361_re <= _T_360_re;
    _T_362_re <= _T_361_re;
    _T_363_re <= _T_362_re;
    _T_364_re <= _T_363_re;
    _T_365_re <= _T_364_re;
    _T_366_re <= _T_365_re;
    _T_367_re <= _T_366_re;
    _T_368_re <= _T_367_re;
    _T_369_re <= _T_368_re;
    _T_370_re <= _T_369_re;
    _T_371_re <= _T_370_re;
    _T_372_re <= _T_371_re;
    _T_373_re <= _T_372_re;
    _T_374_re <= _T_373_re;
    _T_375_re <= _T_374_re;
    _T_376_re <= _T_375_re;
    _T_377_re <= _T_376_re;
    _T_378_re <= _T_377_re;
    _T_379_re <= _T_378_re;
    _T_380_re <= _T_379_re;
    _T_381_re <= _T_380_re;
    _T_382_re <= _T_381_re;
    _T_383_re <= _T_382_re;
    _T_384_re <= _T_383_re;
    _T_385_re <= _T_384_re;
    _T_386_re <= _T_385_re;
    _T_387_re <= _T_386_re;
    _T_388_re <= _T_387_re;
    _T_389_re <= _T_388_re;
    _T_390_re <= _T_389_re;
    _T_391_re <= _T_390_re;
    _T_392_re <= _T_391_re;
    _T_393_re <= _T_392_re;
    _T_394_re <= _T_393_re;
    _T_395_re <= _T_394_re;
    _T_396_re <= _T_395_re;
    _T_397_re <= _T_396_re;
    _T_398_re <= _T_397_re;
    _T_399_re <= _T_398_re;
    _T_400_re <= _T_399_re;
    _T_401_re <= _T_400_re;
    _T_402_re <= _T_401_re;
    _T_403_re <= _T_402_re;
    _T_404_re <= _T_403_re;
    _T_405_re <= _T_404_re;
    _T_406_re <= _T_405_re;
    _T_407_re <= _T_406_re;
    _T_408_re <= _T_407_re;
    _T_410_re <= Butterfly_io_out2_re;
    _T_410_im <= Butterfly_io_out2_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_533_re <= _T_532_re;
    _T_533_im <= _T_532_im;
    _T_534_re <= _T_533_re;
    _T_534_im <= _T_533_im;
    _T_535_re <= _T_534_re;
    _T_535_im <= _T_534_im;
    _T_536_re <= _T_535_re;
    _T_536_im <= _T_535_im;
    _T_537_re <= _T_536_re;
    _T_537_im <= _T_536_im;
    _T_546_re <= Switch_io_out1_re;
    _T_546_im <= Switch_io_out1_im;
    _T_547_re <= _T_546_re;
    _T_547_im <= _T_546_im;
    _T_548_re <= _T_547_re;
    _T_548_im <= _T_547_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_663_re <= _T_662_re;
    _T_663_im <= _T_662_im;
    _T_664_re <= _T_663_re;
    _T_664_im <= _T_663_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_671_re <= _T_670_re;
    _T_671_im <= _T_670_im;
    _T_672_re <= _T_671_re;
    _T_672_im <= _T_671_im;
    _T_673_re <= _T_672_re;
    _T_673_im <= _T_672_im;
    _T_675_re <= Butterfly_1_io_out2_re;
    _T_675_im <= Butterfly_1_io_out2_im;
    _T_676_re <= _T_675_re;
    _T_676_im <= _T_675_im;
    _T_677_re <= _T_676_re;
    _T_677_im <= _T_676_im;
    _T_678_re <= _T_677_re;
    _T_678_im <= _T_677_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_728_re <= _T_727_re;
    _T_728_im <= _T_727_im;
    _T_729_re <= _T_728_re;
    _T_729_im <= _T_728_im;
    _T_730_re <= _T_729_re;
    _T_730_im <= _T_729_im;
    _T_731_re <= _T_730_re;
    _T_731_im <= _T_730_im;
    _T_732_re <= _T_731_re;
    _T_732_im <= _T_731_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_736_re <= _T_735_re;
    _T_736_im <= _T_735_im;
    _T_737_re <= _T_736_re;
    _T_737_im <= _T_736_im;
    _T_738_re <= _T_737_re;
    _T_738_im <= _T_737_im;
    _T_747_re <= Switch_1_io_out1_re;
    _T_747_im <= Switch_1_io_out1_im;
    _T_748_re <= _T_747_re;
    _T_748_im <= _T_747_im;
    _T_749_re <= _T_748_re;
    _T_749_im <= _T_748_im;
    _T_750_re <= _T_749_re;
    _T_750_im <= _T_749_im;
    _T_751_re <= _T_750_re;
    _T_751_im <= _T_750_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_796_re <= _T_795_re;
    _T_796_im <= _T_795_im;
    _T_797_re <= _T_796_re;
    _T_797_im <= _T_796_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_808_re <= _T_807_re;
    _T_808_im <= _T_807_im;
    _T_809_re <= _T_808_re;
    _T_809_im <= _T_808_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_812_re <= Butterfly_2_io_out2_re;
    _T_812_im <= Butterfly_2_io_out2_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_815_re <= _T_814_re;
    _T_815_im <= _T_814_im;
    _T_816_re <= _T_815_re;
    _T_816_im <= _T_815_im;
    _T_817_re <= _T_816_re;
    _T_817_im <= _T_816_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_829_re <= _T_828_re;
    _T_829_im <= _T_828_im;
    _T_830_re <= _T_829_re;
    _T_830_im <= _T_829_im;
    _T_831_re <= _T_830_re;
    _T_831_im <= _T_830_im;
    _T_832_re <= _T_831_re;
    _T_832_im <= _T_831_im;
    _T_833_re <= _T_832_re;
    _T_833_im <= _T_832_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_841_re <= _T_840_re;
    _T_841_im <= _T_840_im;
    _T_842_re <= _T_841_re;
    _T_842_im <= _T_841_im;
    _T_843_re <= _T_842_re;
    _T_843_im <= _T_842_im;
    _T_852_re <= Switch_2_io_out1_re;
    _T_852_im <= Switch_2_io_out1_im;
    _T_853_re <= _T_852_re;
    _T_853_im <= _T_852_im;
    _T_854_re <= _T_853_re;
    _T_854_im <= _T_853_im;
    _T_855_re <= _T_854_re;
    _T_855_im <= _T_854_im;
    _T_856_re <= _T_855_re;
    _T_856_im <= _T_855_im;
    _T_857_re <= _T_856_re;
    _T_857_im <= _T_856_im;
    _T_858_re <= _T_857_re;
    _T_858_im <= _T_857_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_865_re <= _T_864_re;
    _T_865_im <= _T_864_im;
    _T_866_re <= _T_865_re;
    _T_866_im <= _T_865_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_881_re <= _T_880_re;
    _T_881_im <= _T_880_im;
    _T_882_re <= _T_881_re;
    _T_882_im <= _T_881_im;
    _T_883_re <= _T_882_re;
    _T_883_im <= _T_882_im;
    _T_885_re <= Butterfly_3_io_out2_re;
    _T_885_im <= Butterfly_3_io_out2_im;
    _T_886_re <= _T_885_re;
    _T_886_im <= _T_885_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_890_re <= _T_889_re;
    _T_890_im <= _T_889_im;
    _T_891_re <= _T_890_re;
    _T_891_im <= _T_890_im;
    _T_892_re <= _T_891_re;
    _T_892_im <= _T_891_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_898_re <= _T_897_re;
    _T_898_im <= _T_897_im;
    _T_899_re <= _T_898_re;
    _T_899_im <= _T_898_im;
    _T_900_re <= _T_899_re;
    _T_900_im <= _T_899_im;
    _T_909_re <= Switch_3_io_out1_re;
    _T_909_im <= Switch_3_io_out1_im;
    _T_910_re <= _T_909_re;
    _T_910_im <= _T_909_im;
    _T_911_re <= _T_910_re;
    _T_911_im <= _T_910_im;
    _T_912_re <= _T_911_re;
    _T_912_im <= _T_911_im;
    _T_913_re <= _T_912_re;
    _T_913_im <= _T_912_im;
    _T_914_re <= _T_913_re;
    _T_914_im <= _T_913_im;
    _T_915_re <= _T_914_re;
    _T_915_im <= _T_914_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_922_re <= _T_921_re;
    _T_922_im <= _T_921_im;
    _T_923_re <= _T_922_re;
    _T_923_im <= _T_922_im;
    _T_924_re <= _T_923_re;
    _T_924_im <= _T_923_im;
    _T_926_re <= Butterfly_4_io_out2_re;
    _T_926_im <= Butterfly_4_io_out2_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_928_re <= _T_927_re;
    _T_928_im <= _T_927_im;
    _T_929_re <= _T_928_re;
    _T_929_im <= _T_928_im;
    _T_930_re <= _T_929_re;
    _T_930_im <= _T_929_im;
    _T_931_re <= _T_930_re;
    _T_931_im <= _T_930_im;
    _T_932_re <= _T_931_re;
    _T_932_im <= _T_931_im;
    _T_933_re <= _T_932_re;
    _T_933_im <= _T_932_im;
    _T_942_re <= Switch_4_io_out1_re;
    _T_942_im <= Switch_4_io_out1_im;
    _T_943_re <= _T_942_re;
    _T_943_im <= _T_942_im;
    _T_944_re <= _T_943_re;
    _T_944_im <= _T_943_im;
    _T_945_re <= _T_944_re;
    _T_945_im <= _T_944_im;
    _T_946_re <= _T_945_re;
    _T_946_im <= _T_945_im;
    _T_947_re <= _T_946_re;
    _T_947_im <= _T_946_im;
    _T_948_re <= _T_947_re;
    _T_948_im <= _T_947_im;
    _T_949_re <= _T_948_re;
    _T_949_im <= _T_948_im;
    _T_951_re <= Butterfly_5_io_out2_re;
    _T_951_im <= Butterfly_5_io_out2_im;
    _T_952_re <= _T_951_re;
    _T_952_im <= _T_951_im;
    _T_953_re <= _T_952_re;
    _T_953_im <= _T_952_im;
    _T_954_re <= _T_953_re;
    _T_954_im <= _T_953_im;
    _T_963_re <= Switch_5_io_out1_re;
    _T_963_im <= Switch_5_io_out1_im;
    _T_964_re <= _T_963_re;
    _T_964_im <= _T_963_im;
    _T_965_re <= _T_964_re;
    _T_965_im <= _T_964_im;
    _T_966_re <= _T_965_re;
    _T_966_im <= _T_965_im;
    _T_968_re <= Butterfly_6_io_out2_re;
    _T_968_im <= Butterfly_6_io_out2_im;
    _T_969_re <= _T_968_re;
    _T_969_im <= _T_968_im;
    _T_978_re <= Switch_6_io_out1_re;
    _T_978_im <= Switch_6_io_out1_im;
    _T_979_re <= _T_978_re;
    _T_979_im <= _T_978_im;
    _T_981_re <= Butterfly_7_io_out2_re;
    _T_981_im <= Butterfly_7_io_out2_im;
    out1D1_re <= Switch_7_io_out1_re;
    out1D1_im <= Switch_7_io_out1_im;
    _T_988_re <= ComplexAdd_io_res_re;
    _T_988_im <= ComplexAdd_io_res_im;
    _T_989_re <= ComplexSub_io_res_re;
    _T_989_im <= ComplexSub_io_res_im;
    _T_990 <= cnt;
  end
endmodule
module Reorder(
  input         clock,
  input         reset,
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_in_valid,
  output [31:0] io_out_re,
  output [31:0] io_out_im,
  output        io_out_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rambank0_re [0:255]; // @[Reorder.scala 18:21]
  wire [31:0] rambank0_re__T_80_data; // @[Reorder.scala 18:21]
  wire [7:0] rambank0_re__T_80_addr; // @[Reorder.scala 18:21]
  wire [31:0] rambank0_re__T_69_data; // @[Reorder.scala 18:21]
  wire [7:0] rambank0_re__T_69_addr; // @[Reorder.scala 18:21]
  wire  rambank0_re__T_69_mask; // @[Reorder.scala 18:21]
  wire  rambank0_re__T_69_en; // @[Reorder.scala 18:21]
  reg [31:0] rambank0_im [0:255]; // @[Reorder.scala 18:21]
  wire [31:0] rambank0_im__T_80_data; // @[Reorder.scala 18:21]
  wire [7:0] rambank0_im__T_80_addr; // @[Reorder.scala 18:21]
  wire [31:0] rambank0_im__T_69_data; // @[Reorder.scala 18:21]
  wire [7:0] rambank0_im__T_69_addr; // @[Reorder.scala 18:21]
  wire  rambank0_im__T_69_mask; // @[Reorder.scala 18:21]
  wire  rambank0_im__T_69_en; // @[Reorder.scala 18:21]
  reg [31:0] rambank1_re [0:255]; // @[Reorder.scala 19:21]
  wire [31:0] rambank1_re__T_82_data; // @[Reorder.scala 19:21]
  wire [7:0] rambank1_re__T_82_addr; // @[Reorder.scala 19:21]
  wire [31:0] rambank1_re__T_71_data; // @[Reorder.scala 19:21]
  wire [7:0] rambank1_re__T_71_addr; // @[Reorder.scala 19:21]
  wire  rambank1_re__T_71_mask; // @[Reorder.scala 19:21]
  wire  rambank1_re__T_71_en; // @[Reorder.scala 19:21]
  reg [31:0] rambank1_im [0:255]; // @[Reorder.scala 19:21]
  wire [31:0] rambank1_im__T_82_data; // @[Reorder.scala 19:21]
  wire [7:0] rambank1_im__T_82_addr; // @[Reorder.scala 19:21]
  wire [31:0] rambank1_im__T_71_data; // @[Reorder.scala 19:21]
  wire [7:0] rambank1_im__T_71_addr; // @[Reorder.scala 19:21]
  wire  rambank1_im__T_71_mask; // @[Reorder.scala 19:21]
  wire  rambank1_im__T_71_en; // @[Reorder.scala 19:21]
  reg [7:0] in_counter; // @[Reorder.scala 22:27]
  reg [8:0] out_counter; // @[Reorder.scala 23:28]
  wire [8:0] _T = {in_counter,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_5 = {{4'd0}, _T[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_7 = {_T[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_9 = _T_7 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_10 = _T_5 | _T_9; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_19 = {{2'd0}, _T_10[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_15 = _GEN_19 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_17 = {_T_10[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_19 = _T_17 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_20 = _T_15 | _T_19; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_20 = {{1'd0}, _T_20[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_25 = _GEN_20 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_27 = {_T_20[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_29 = _T_27 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_30 = _T_25 | _T_29; // @[Bitwise.scala 103:39]
  wire [8:0] index1 = {_T_30,_T[8]}; // @[Cat.scala 29:58]
  wire [8:0] _T_32 = {in_counter,1'h1}; // @[Cat.scala 29:58]
  wire [7:0] _T_37 = {{4'd0}, _T_32[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_39 = {_T_32[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_41 = _T_39 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_21 = {{2'd0}, _T_42[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_47 = _GEN_21 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_49 = {_T_42[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_51 = _T_49 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_22 = {{1'd0}, _T_52[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_57 = _GEN_22 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_59 = {_T_52[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_61 = _T_59 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39]
  wire [8:0] index2 = {_T_62,_T_32[8]}; // @[Cat.scala 29:58]
  wire  _T_64 = in_counter != 8'h0; // @[Reorder.scala 26:34]
  wire  _T_65 = io_in_valid | _T_64; // @[Reorder.scala 26:20]
  wire [7:0] _T_67 = in_counter + 8'h1; // @[Reorder.scala 27:30]
  reg [7:0] _T_72; // @[Reorder.scala 32:27]
  wire  _T_73 = _T_72 == 8'hff; // @[Reorder.scala 32:40]
  wire  _T_74 = out_counter != 9'h0; // @[Reorder.scala 32:90]
  wire [8:0] _T_77 = out_counter + 9'h1; // @[Reorder.scala 34:32]
  wire  _T_78 = out_counter < 9'h100; // @[Reorder.scala 37:20]
  assign rambank0_re__T_80_addr = out_counter[7:0];
  assign rambank0_re__T_80_data = rambank0_re[rambank0_re__T_80_addr]; // @[Reorder.scala 18:21]
  assign rambank0_re__T_69_data = io_in1_re;
  assign rambank0_re__T_69_addr = index1[7:0];
  assign rambank0_re__T_69_mask = 1'h1;
  assign rambank0_re__T_69_en = io_in_valid | _T_64;
  assign rambank0_im__T_80_addr = out_counter[7:0];
  assign rambank0_im__T_80_data = rambank0_im[rambank0_im__T_80_addr]; // @[Reorder.scala 18:21]
  assign rambank0_im__T_69_data = io_in1_im;
  assign rambank0_im__T_69_addr = index1[7:0];
  assign rambank0_im__T_69_mask = 1'h1;
  assign rambank0_im__T_69_en = io_in_valid | _T_64;
  assign rambank1_re__T_82_addr = out_counter[7:0];
  assign rambank1_re__T_82_data = rambank1_re[rambank1_re__T_82_addr]; // @[Reorder.scala 19:21]
  assign rambank1_re__T_71_data = io_in2_re;
  assign rambank1_re__T_71_addr = index2[7:0];
  assign rambank1_re__T_71_mask = 1'h1;
  assign rambank1_re__T_71_en = io_in_valid | _T_64;
  assign rambank1_im__T_82_addr = out_counter[7:0];
  assign rambank1_im__T_82_data = rambank1_im[rambank1_im__T_82_addr]; // @[Reorder.scala 19:21]
  assign rambank1_im__T_71_data = io_in2_im;
  assign rambank1_im__T_71_addr = index2[7:0];
  assign rambank1_im__T_71_mask = 1'h1;
  assign rambank1_im__T_71_en = io_in_valid | _T_64;
  assign io_out_re = _T_78 ? $signed(rambank0_re__T_80_data) : $signed(rambank1_re__T_82_data); // @[Reorder.scala 38:12 Reorder.scala 40:12]
  assign io_out_im = _T_78 ? $signed(rambank0_im__T_80_data) : $signed(rambank1_im__T_82_data); // @[Reorder.scala 38:12 Reorder.scala 40:12]
  assign io_out_valid = _T_73 | _T_74; // @[Reorder.scala 32:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank0_re[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank0_im[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank1_re[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank1_im[initvar] = _RAND_3[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_counter = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  out_counter = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  _T_72 = _RAND_6[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(rambank0_re__T_69_en & rambank0_re__T_69_mask) begin
      rambank0_re[rambank0_re__T_69_addr] <= rambank0_re__T_69_data; // @[Reorder.scala 18:21]
    end
    if(rambank0_im__T_69_en & rambank0_im__T_69_mask) begin
      rambank0_im[rambank0_im__T_69_addr] <= rambank0_im__T_69_data; // @[Reorder.scala 18:21]
    end
    if(rambank1_re__T_71_en & rambank1_re__T_71_mask) begin
      rambank1_re[rambank1_re__T_71_addr] <= rambank1_re__T_71_data; // @[Reorder.scala 19:21]
    end
    if(rambank1_im__T_71_en & rambank1_im__T_71_mask) begin
      rambank1_im[rambank1_im__T_71_addr] <= rambank1_im__T_71_data; // @[Reorder.scala 19:21]
    end
    if (reset) begin
      in_counter <= 8'h0;
    end else if (_T_65) begin
      in_counter <= _T_67;
    end
    if (reset) begin
      out_counter <= 9'h0;
    end else if (io_out_valid) begin
      out_counter <= _T_77;
    end
    _T_72 <= in_counter;
  end
endmodule
module FFTReorder(
  input         clock,
  input         reset,
  input  [31:0] io_dIn_re,
  input         io_din_valid,
  output [31:0] io_dOut_re,
  output [31:0] io_dOut_im,
  output        io_dout_valid,
  output        io_busy
);
  wire  fftblock_clock; // @[Reorder.scala 56:29]
  wire  fftblock_reset; // @[Reorder.scala 56:29]
  wire [31:0] fftblock_io_dIn_re; // @[Reorder.scala 56:29]
  wire  fftblock_io_din_valid; // @[Reorder.scala 56:29]
  wire [31:0] fftblock_io_dOut1_re; // @[Reorder.scala 56:29]
  wire [31:0] fftblock_io_dOut1_im; // @[Reorder.scala 56:29]
  wire [31:0] fftblock_io_dOut2_re; // @[Reorder.scala 56:29]
  wire [31:0] fftblock_io_dOut2_im; // @[Reorder.scala 56:29]
  wire  fftblock_io_dout_valid; // @[Reorder.scala 56:29]
  wire  fftblock_io_busy; // @[Reorder.scala 56:29]
  wire  reorderblock_clock; // @[Reorder.scala 60:28]
  wire  reorderblock_reset; // @[Reorder.scala 60:28]
  wire [31:0] reorderblock_io_in1_re; // @[Reorder.scala 60:28]
  wire [31:0] reorderblock_io_in1_im; // @[Reorder.scala 60:28]
  wire [31:0] reorderblock_io_in2_re; // @[Reorder.scala 60:28]
  wire [31:0] reorderblock_io_in2_im; // @[Reorder.scala 60:28]
  wire  reorderblock_io_in_valid; // @[Reorder.scala 60:28]
  wire [31:0] reorderblock_io_out_re; // @[Reorder.scala 60:28]
  wire [31:0] reorderblock_io_out_im; // @[Reorder.scala 60:28]
  wire  reorderblock_io_out_valid; // @[Reorder.scala 60:28]
  FFT fftblock ( // @[Reorder.scala 56:29]
    .clock(fftblock_clock),
    .reset(fftblock_reset),
    .io_dIn_re(fftblock_io_dIn_re),
    .io_din_valid(fftblock_io_din_valid),
    .io_dOut1_re(fftblock_io_dOut1_re),
    .io_dOut1_im(fftblock_io_dOut1_im),
    .io_dOut2_re(fftblock_io_dOut2_re),
    .io_dOut2_im(fftblock_io_dOut2_im),
    .io_dout_valid(fftblock_io_dout_valid),
    .io_busy(fftblock_io_busy)
  );
  Reorder reorderblock ( // @[Reorder.scala 60:28]
    .clock(reorderblock_clock),
    .reset(reorderblock_reset),
    .io_in1_re(reorderblock_io_in1_re),
    .io_in1_im(reorderblock_io_in1_im),
    .io_in2_re(reorderblock_io_in2_re),
    .io_in2_im(reorderblock_io_in2_im),
    .io_in_valid(reorderblock_io_in_valid),
    .io_out_re(reorderblock_io_out_re),
    .io_out_im(reorderblock_io_out_im),
    .io_out_valid(reorderblock_io_out_valid)
  );
  assign io_dOut_re = reorderblock_io_out_re; // @[Reorder.scala 65:11]
  assign io_dOut_im = reorderblock_io_out_im; // @[Reorder.scala 65:11]
  assign io_dout_valid = reorderblock_io_out_valid; // @[Reorder.scala 66:17]
  assign io_busy = fftblock_io_busy; // @[Reorder.scala 67:11]
  assign fftblock_clock = clock;
  assign fftblock_reset = reset;
  assign fftblock_io_dIn_re = io_dIn_re; // @[Reorder.scala 57:19]
  assign fftblock_io_din_valid = io_din_valid; // @[Reorder.scala 58:25]
  assign reorderblock_clock = clock;
  assign reorderblock_reset = reset;
  assign reorderblock_io_in1_re = fftblock_io_dOut1_re; // @[Reorder.scala 61:23]
  assign reorderblock_io_in1_im = fftblock_io_dOut1_im; // @[Reorder.scala 61:23]
  assign reorderblock_io_in2_re = fftblock_io_dOut2_re; // @[Reorder.scala 62:23]
  assign reorderblock_io_in2_im = fftblock_io_dOut2_im; // @[Reorder.scala 62:23]
  assign reorderblock_io_in_valid = fftblock_io_dout_valid; // @[Reorder.scala 63:28]
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_re,
  input  [31:0] io_enq_bits_im,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_re,
  output [31:0] io_deq_bits_im
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_re [0:1023]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_re__T_15_data; // @[Decoupled.scala 209:16]
  wire [9:0] ram_re__T_15_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_re__T_5_data; // @[Decoupled.scala 209:16]
  wire [9:0] ram_re__T_5_addr; // @[Decoupled.scala 209:16]
  wire  ram_re__T_5_mask; // @[Decoupled.scala 209:16]
  wire  ram_re__T_5_en; // @[Decoupled.scala 209:16]
  reg [31:0] ram_im [0:1023]; // @[Decoupled.scala 209:16]
  wire [31:0] ram_im__T_15_data; // @[Decoupled.scala 209:16]
  wire [9:0] ram_im__T_15_addr; // @[Decoupled.scala 209:16]
  wire [31:0] ram_im__T_5_data; // @[Decoupled.scala 209:16]
  wire [9:0] ram_im__T_5_addr; // @[Decoupled.scala 209:16]
  wire  ram_im__T_5_mask; // @[Decoupled.scala 209:16]
  wire  ram_im__T_5_en; // @[Decoupled.scala 209:16]
  reg [9:0] _T; // @[Counter.scala 29:33]
  reg [9:0] _T_1; // @[Counter.scala 29:33]
  reg  maybe_full; // @[Decoupled.scala 212:27]
  wire  ptr_match = _T == _T_1; // @[Decoupled.scala 214:33]
  wire  _T_2 = ~maybe_full; // @[Decoupled.scala 215:28]
  wire  empty = ptr_match & _T_2; // @[Decoupled.scala 215:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 216:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [9:0] _T_8 = _T + 10'h1; // @[Counter.scala 39:22]
  wire [9:0] _T_11 = _T_1 + 10'h1; // @[Counter.scala 39:22]
  wire  _T_12 = do_enq != do_deq; // @[Decoupled.scala 227:16]
  assign ram_re__T_15_addr = _T_1;
  assign ram_re__T_15_data = ram_re[ram_re__T_15_addr]; // @[Decoupled.scala 209:16]
  assign ram_re__T_5_data = io_enq_bits_re;
  assign ram_re__T_5_addr = _T;
  assign ram_re__T_5_mask = 1'h1;
  assign ram_re__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_im__T_15_addr = _T_1;
  assign ram_im__T_15_data = ram_im[ram_im__T_15_addr]; // @[Decoupled.scala 209:16]
  assign ram_im__T_5_data = io_enq_bits_im;
  assign ram_im__T_5_addr = _T;
  assign ram_im__T_5_mask = 1'h1;
  assign ram_im__T_5_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 231:16]
  assign io_deq_bits_re = ram_re__T_15_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_im = ram_im__T_15_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram_re[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram_im[initvar] = _RAND_1[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_re__T_5_en & ram_re__T_5_mask) begin
      ram_re[ram_re__T_5_addr] <= ram_re__T_5_data; // @[Decoupled.scala 209:16]
    end
    if(ram_im__T_5_en & ram_im__T_5_mask) begin
      ram_im[ram_im__T_5_addr] <= ram_im__T_5_data; // @[Decoupled.scala 209:16]
    end
    if (reset) begin
      _T <= 10'h0;
    end else if (do_enq) begin
      _T <= _T_8;
    end
    if (reset) begin
      _T_1 <= 10'h0;
    end else if (do_deq) begin
      _T_1 <= _T_11;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module TOP(
  input         clock,
  input         reset,
  output        io_din_ready,
  input         io_din_valid,
  input  [31:0] io_din_bits_re,
  input         io_dout_ready,
  output        io_dout_valid,
  output [31:0] io_dout_bits_re,
  output [31:0] io_dout_bits_im
);
  wire  FFT_clock; // @[TOP.scala 21:19]
  wire  FFT_reset; // @[TOP.scala 21:19]
  wire [31:0] FFT_io_dIn_re; // @[TOP.scala 21:19]
  wire  FFT_io_din_valid; // @[TOP.scala 21:19]
  wire [31:0] FFT_io_dOut_re; // @[TOP.scala 21:19]
  wire [31:0] FFT_io_dOut_im; // @[TOP.scala 21:19]
  wire  FFT_io_dout_valid; // @[TOP.scala 21:19]
  wire  FFT_io_busy; // @[TOP.scala 21:19]
  wire  FIFO_clock; // @[Decoupled.scala 287:21]
  wire  FIFO_reset; // @[Decoupled.scala 287:21]
  wire  FIFO_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  FIFO_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] FIFO_io_enq_bits_re; // @[Decoupled.scala 287:21]
  wire [31:0] FIFO_io_enq_bits_im; // @[Decoupled.scala 287:21]
  wire  FIFO_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  FIFO_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] FIFO_io_deq_bits_re; // @[Decoupled.scala 287:21]
  wire [31:0] FIFO_io_deq_bits_im; // @[Decoupled.scala 287:21]
  wire  _T = ~FFT_io_busy; // @[TOP.scala 28:36]
  wire  FIFOcmd_ready = FIFO_io_enq_ready; // @[TOP.scala 22:21 Decoupled.scala 290:17]
  FFTReorder FFT ( // @[TOP.scala 21:19]
    .clock(FFT_clock),
    .reset(FFT_reset),
    .io_dIn_re(FFT_io_dIn_re),
    .io_din_valid(FFT_io_din_valid),
    .io_dOut_re(FFT_io_dOut_re),
    .io_dOut_im(FFT_io_dOut_im),
    .io_dout_valid(FFT_io_dout_valid),
    .io_busy(FFT_io_busy)
  );
  Queue FIFO ( // @[Decoupled.scala 287:21]
    .clock(FIFO_clock),
    .reset(FIFO_reset),
    .io_enq_ready(FIFO_io_enq_ready),
    .io_enq_valid(FIFO_io_enq_valid),
    .io_enq_bits_re(FIFO_io_enq_bits_re),
    .io_enq_bits_im(FIFO_io_enq_bits_im),
    .io_deq_ready(FIFO_io_deq_ready),
    .io_deq_valid(FIFO_io_deq_valid),
    .io_deq_bits_re(FIFO_io_deq_bits_re),
    .io_deq_bits_im(FIFO_io_deq_bits_im)
  );
  assign io_din_ready = FIFOcmd_ready & _T; // @[TOP.scala 28:16]
  assign io_dout_valid = FIFO_io_deq_ready & FIFO_io_deq_valid; // @[TOP.scala 32:17]
  assign io_dout_bits_re = FIFO_io_deq_bits_re; // @[TOP.scala 33:16]
  assign io_dout_bits_im = FIFO_io_deq_bits_im; // @[TOP.scala 33:16]
  assign FFT_clock = clock;
  assign FFT_reset = reset;
  assign FFT_io_dIn_re = io_din_bits_re; // @[TOP.scala 30:14]
  assign FFT_io_din_valid = io_din_ready & io_din_valid; // @[TOP.scala 29:20]
  assign FIFO_clock = clock;
  assign FIFO_reset = reset;
  assign FIFO_io_enq_valid = FFT_io_dout_valid; // @[Decoupled.scala 288:22]
  assign FIFO_io_enq_bits_re = FFT_io_dOut_re; // @[Decoupled.scala 289:21]
  assign FIFO_io_enq_bits_im = FFT_io_dOut_im; // @[Decoupled.scala 289:21]
  assign FIFO_io_deq_ready = io_dout_ready; // @[TOP.scala 26:14]
endmodule
module ComplexEnergy(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_value
);
  wire [63:0] _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 61:29]
  wire [63:0] _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 61:53]
  wire [63:0] _T_4 = $signed(_T) + $signed(_T_1); // @[Butterfly.scala 61:41]
  wire [47:0] _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 61:16]
  assign io_res_value = _GEN_0[31:0]; // @[Butterfly.scala 61:16]
endmodule
module SpectrogramGen(
  input         clock,
  input         reset,
  output        io_FFTsignal_ready,
  input         io_FFTsignal_valid,
  input  [31:0] io_FFTsignal_bits_re,
  input  [31:0] io_FFTsignal_bits_im,
  input         io_Spectrogram_ready,
  output        io_Spectrogram_valid,
  output [31:0] io_Spectrogram_bits_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] ComplexEnergy_io_op1_re; // @[Butterfly.scala 65:22]
  wire [31:0] ComplexEnergy_io_op1_im; // @[Butterfly.scala 65:22]
  wire [31:0] ComplexEnergy_io_op2_re; // @[Butterfly.scala 65:22]
  wire [31:0] ComplexEnergy_io_op2_im; // @[Butterfly.scala 65:22]
  wire [31:0] ComplexEnergy_io_res_value; // @[Butterfly.scala 65:22]
  reg [31:0] SpectrogramReg_value; // @[SpectrogramGen.scala 18:27]
  reg [9:0] SpectrogramCnt; // @[SpectrogramGen.scala 19:31]
  reg  Spectrogram_valid; // @[SpectrogramGen.scala 20:34]
  wire  _T = io_FFTsignal_valid & io_Spectrogram_ready; // @[SpectrogramGen.scala 22:28]
  wire  _T_1 = SpectrogramCnt < 10'h101; // @[SpectrogramGen.scala 24:25]
  wire [9:0] _T_3 = SpectrogramCnt + 10'h1; // @[SpectrogramGen.scala 26:40]
  wire  _T_4 = SpectrogramCnt < 10'h200; // @[SpectrogramGen.scala 27:31]
  ComplexEnergy ComplexEnergy ( // @[Butterfly.scala 65:22]
    .io_op1_re(ComplexEnergy_io_op1_re),
    .io_op1_im(ComplexEnergy_io_op1_im),
    .io_op2_re(ComplexEnergy_io_op2_re),
    .io_op2_im(ComplexEnergy_io_op2_im),
    .io_res_value(ComplexEnergy_io_res_value)
  );
  assign io_FFTsignal_ready = io_Spectrogram_ready; // @[SpectrogramGen.scala 48:22]
  assign io_Spectrogram_valid = Spectrogram_valid; // @[SpectrogramGen.scala 50:24]
  assign io_Spectrogram_bits_value = SpectrogramReg_value; // @[SpectrogramGen.scala 49:23]
  assign ComplexEnergy_io_op1_re = io_FFTsignal_bits_re; // @[Butterfly.scala 66:17]
  assign ComplexEnergy_io_op1_im = io_FFTsignal_bits_im; // @[Butterfly.scala 66:17]
  assign ComplexEnergy_io_op2_re = io_FFTsignal_bits_re; // @[Butterfly.scala 67:17]
  assign ComplexEnergy_io_op2_im = io_FFTsignal_bits_im; // @[Butterfly.scala 67:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  SpectrogramReg_value = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  SpectrogramCnt = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  Spectrogram_valid = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      SpectrogramReg_value <= ComplexEnergy_io_res_value;
    end
    if (reset) begin
      SpectrogramCnt <= 10'h0;
    end else if (_T) begin
      if (_T_1) begin
        SpectrogramCnt <= _T_3;
      end else if (_T_4) begin
        SpectrogramCnt <= _T_3;
      end else begin
        SpectrogramCnt <= 10'h0;
      end
    end
    if (reset) begin
      Spectrogram_valid <= 1'h0;
    end else if (_T) begin
      Spectrogram_valid <= _T_1;
    end
  end
endmodule
module SpectrogramGenWithFIFO(
  input         clock,
  input         reset,
  output        io_FFTsignal_ready,
  input         io_FFTsignal_valid,
  input  [31:0] io_FFTsignal_bits_re,
  input  [31:0] io_FFTsignal_bits_im,
  input         io_Spectrogram_ready,
  output        io_Spectrogram_valid,
  output [31:0] io_Spectrogram_bits_value
);
  wire  SpectrogramGenblock_clock; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire  SpectrogramGenblock_reset; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire  SpectrogramGenblock_io_FFTsignal_ready; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire  SpectrogramGenblock_io_FFTsignal_valid; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire [31:0] SpectrogramGenblock_io_FFTsignal_bits_re; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire [31:0] SpectrogramGenblock_io_FFTsignal_bits_im; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire  SpectrogramGenblock_io_Spectrogram_ready; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire  SpectrogramGenblock_io_Spectrogram_valid; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire [31:0] SpectrogramGenblock_io_Spectrogram_bits_value; // @[SpectrogramGenWithFIFO.scala 17:51]
  wire  SpectrogramFIFO_clock; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire  SpectrogramFIFO_reset; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire [31:0] SpectrogramFIFO_io_datain_value; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire [31:0] SpectrogramFIFO_io_dataout_value; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire  SpectrogramFIFO_io_wr; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire  SpectrogramFIFO_io_rd; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire  SpectrogramFIFO_io_full; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire  SpectrogramFIFO_io_empty; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire  SpectrogramFIFO_io_MorethanN; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire [31:0] SpectrogramFIFO_io_count; // @[SpectrogramGenWithFIFO.scala 18:39]
  wire [31:0] _T_1 = 32'h400 - SpectrogramFIFO_io_count; // @[SpectrogramGenWithFIFO.scala 23:67]
  wire  _T_4 = ~SpectrogramFIFO_io_empty; // @[SpectrogramGenWithFIFO.scala 27:33]
  wire  _T_5 = SpectrogramFIFO_io_wr & SpectrogramFIFO_io_empty; // @[SpectrogramGenWithFIFO.scala 27:85]
  SpectrogramGen SpectrogramGenblock ( // @[SpectrogramGenWithFIFO.scala 17:51]
    .clock(SpectrogramGenblock_clock),
    .reset(SpectrogramGenblock_reset),
    .io_FFTsignal_ready(SpectrogramGenblock_io_FFTsignal_ready),
    .io_FFTsignal_valid(SpectrogramGenblock_io_FFTsignal_valid),
    .io_FFTsignal_bits_re(SpectrogramGenblock_io_FFTsignal_bits_re),
    .io_FFTsignal_bits_im(SpectrogramGenblock_io_FFTsignal_bits_im),
    .io_Spectrogram_ready(SpectrogramGenblock_io_Spectrogram_ready),
    .io_Spectrogram_valid(SpectrogramGenblock_io_Spectrogram_valid),
    .io_Spectrogram_bits_value(SpectrogramGenblock_io_Spectrogram_bits_value)
  );
  MyFifo SpectrogramFIFO ( // @[SpectrogramGenWithFIFO.scala 18:39]
    .clock(SpectrogramFIFO_clock),
    .reset(SpectrogramFIFO_reset),
    .io_datain_value(SpectrogramFIFO_io_datain_value),
    .io_dataout_value(SpectrogramFIFO_io_dataout_value),
    .io_wr(SpectrogramFIFO_io_wr),
    .io_rd(SpectrogramFIFO_io_rd),
    .io_full(SpectrogramFIFO_io_full),
    .io_empty(SpectrogramFIFO_io_empty),
    .io_MorethanN(SpectrogramFIFO_io_MorethanN),
    .io_count(SpectrogramFIFO_io_count)
  );
  assign io_FFTsignal_ready = SpectrogramGenblock_io_FFTsignal_ready; // @[SpectrogramGenWithFIFO.scala 20:16]
  assign io_Spectrogram_valid = _T_4 | _T_5; // @[SpectrogramGenWithFIFO.scala 27:30]
  assign io_Spectrogram_bits_value = SpectrogramFIFO_io_dataout_value; // @[SpectrogramGenWithFIFO.scala 28:30]
  assign SpectrogramGenblock_clock = clock;
  assign SpectrogramGenblock_reset = reset;
  assign SpectrogramGenblock_io_FFTsignal_valid = io_FFTsignal_valid; // @[SpectrogramGenWithFIFO.scala 20:16]
  assign SpectrogramGenblock_io_FFTsignal_bits_re = io_FFTsignal_bits_re; // @[SpectrogramGenWithFIFO.scala 20:16]
  assign SpectrogramGenblock_io_FFTsignal_bits_im = io_FFTsignal_bits_im; // @[SpectrogramGenWithFIFO.scala 20:16]
  assign SpectrogramGenblock_io_Spectrogram_ready = _T_1 > 32'h101; // @[SpectrogramGenWithFIFO.scala 23:44]
  assign SpectrogramFIFO_clock = clock;
  assign SpectrogramFIFO_reset = reset;
  assign SpectrogramFIFO_io_datain_value = SpectrogramGenblock_io_Spectrogram_bits_value; // @[SpectrogramGenWithFIFO.scala 24:30]
  assign SpectrogramFIFO_io_wr = SpectrogramGenblock_io_Spectrogram_valid; // @[SpectrogramGenWithFIFO.scala 25:30]
  assign SpectrogramFIFO_io_rd = io_Spectrogram_ready & io_Spectrogram_valid; // @[SpectrogramGenWithFIFO.scala 26:30]
endmodule
module STFT(
  input         clock,
  input         reset,
  output        io_signal_ready,
  input         io_signal_valid,
  input  [31:0] io_signal_bits_value,
  output        io_cosines_ready,
  input         io_cosines_valid,
  input  [31:0] io_cosines_bits_value,
  input         io_spectrogram_ready,
  output        io_spectrogram_valid,
  output [31:0] io_spectrogram_bits_value
);
  wire  HanningBlock_clock; // @[STFT.scala 26:45]
  wire  HanningBlock_reset; // @[STFT.scala 26:45]
  wire  HanningBlock_io_signal_ready; // @[STFT.scala 26:45]
  wire  HanningBlock_io_signal_valid; // @[STFT.scala 26:45]
  wire [31:0] HanningBlock_io_signal_bits_value; // @[STFT.scala 26:45]
  wire  HanningBlock_io_cosines_ready; // @[STFT.scala 26:45]
  wire  HanningBlock_io_cosines_valid; // @[STFT.scala 26:45]
  wire [31:0] HanningBlock_io_cosines_bits_value; // @[STFT.scala 26:45]
  wire  HanningBlock_io_HanningSignal_ready; // @[STFT.scala 26:45]
  wire  HanningBlock_io_HanningSignal_valid; // @[STFT.scala 26:45]
  wire [31:0] HanningBlock_io_HanningSignal_bits_value; // @[STFT.scala 26:45]
  wire  FFTBlock_clock; // @[STFT.scala 27:29]
  wire  FFTBlock_reset; // @[STFT.scala 27:29]
  wire  FFTBlock_io_din_ready; // @[STFT.scala 27:29]
  wire  FFTBlock_io_din_valid; // @[STFT.scala 27:29]
  wire [31:0] FFTBlock_io_din_bits_re; // @[STFT.scala 27:29]
  wire  FFTBlock_io_dout_ready; // @[STFT.scala 27:29]
  wire  FFTBlock_io_dout_valid; // @[STFT.scala 27:29]
  wire [31:0] FFTBlock_io_dout_bits_re; // @[STFT.scala 27:29]
  wire [31:0] FFTBlock_io_dout_bits_im; // @[STFT.scala 27:29]
  wire  SpectrogramGenBlock_clock; // @[STFT.scala 28:59]
  wire  SpectrogramGenBlock_reset; // @[STFT.scala 28:59]
  wire  SpectrogramGenBlock_io_FFTsignal_ready; // @[STFT.scala 28:59]
  wire  SpectrogramGenBlock_io_FFTsignal_valid; // @[STFT.scala 28:59]
  wire [31:0] SpectrogramGenBlock_io_FFTsignal_bits_re; // @[STFT.scala 28:59]
  wire [31:0] SpectrogramGenBlock_io_FFTsignal_bits_im; // @[STFT.scala 28:59]
  wire  SpectrogramGenBlock_io_Spectrogram_ready; // @[STFT.scala 28:59]
  wire  SpectrogramGenBlock_io_Spectrogram_valid; // @[STFT.scala 28:59]
  wire [31:0] SpectrogramGenBlock_io_Spectrogram_bits_value; // @[STFT.scala 28:59]
  HanningWithFIFO HanningBlock ( // @[STFT.scala 26:45]
    .clock(HanningBlock_clock),
    .reset(HanningBlock_reset),
    .io_signal_ready(HanningBlock_io_signal_ready),
    .io_signal_valid(HanningBlock_io_signal_valid),
    .io_signal_bits_value(HanningBlock_io_signal_bits_value),
    .io_cosines_ready(HanningBlock_io_cosines_ready),
    .io_cosines_valid(HanningBlock_io_cosines_valid),
    .io_cosines_bits_value(HanningBlock_io_cosines_bits_value),
    .io_HanningSignal_ready(HanningBlock_io_HanningSignal_ready),
    .io_HanningSignal_valid(HanningBlock_io_HanningSignal_valid),
    .io_HanningSignal_bits_value(HanningBlock_io_HanningSignal_bits_value)
  );
  TOP FFTBlock ( // @[STFT.scala 27:29]
    .clock(FFTBlock_clock),
    .reset(FFTBlock_reset),
    .io_din_ready(FFTBlock_io_din_ready),
    .io_din_valid(FFTBlock_io_din_valid),
    .io_din_bits_re(FFTBlock_io_din_bits_re),
    .io_dout_ready(FFTBlock_io_dout_ready),
    .io_dout_valid(FFTBlock_io_dout_valid),
    .io_dout_bits_re(FFTBlock_io_dout_bits_re),
    .io_dout_bits_im(FFTBlock_io_dout_bits_im)
  );
  SpectrogramGenWithFIFO SpectrogramGenBlock ( // @[STFT.scala 28:59]
    .clock(SpectrogramGenBlock_clock),
    .reset(SpectrogramGenBlock_reset),
    .io_FFTsignal_ready(SpectrogramGenBlock_io_FFTsignal_ready),
    .io_FFTsignal_valid(SpectrogramGenBlock_io_FFTsignal_valid),
    .io_FFTsignal_bits_re(SpectrogramGenBlock_io_FFTsignal_bits_re),
    .io_FFTsignal_bits_im(SpectrogramGenBlock_io_FFTsignal_bits_im),
    .io_Spectrogram_ready(SpectrogramGenBlock_io_Spectrogram_ready),
    .io_Spectrogram_valid(SpectrogramGenBlock_io_Spectrogram_valid),
    .io_Spectrogram_bits_value(SpectrogramGenBlock_io_Spectrogram_bits_value)
  );
  assign io_signal_ready = HanningBlock_io_signal_ready; // @[STFT.scala 30:13]
  assign io_cosines_ready = HanningBlock_io_cosines_ready; // @[STFT.scala 31:14]
  assign io_spectrogram_valid = SpectrogramGenBlock_io_Spectrogram_valid; // @[STFT.scala 39:18]
  assign io_spectrogram_bits_value = SpectrogramGenBlock_io_Spectrogram_bits_value; // @[STFT.scala 39:18]
  assign HanningBlock_clock = clock;
  assign HanningBlock_reset = reset;
  assign HanningBlock_io_signal_valid = io_signal_valid; // @[STFT.scala 30:13]
  assign HanningBlock_io_signal_bits_value = io_signal_bits_value; // @[STFT.scala 30:13]
  assign HanningBlock_io_cosines_valid = io_cosines_valid; // @[STFT.scala 31:14]
  assign HanningBlock_io_cosines_bits_value = io_cosines_bits_value; // @[STFT.scala 31:14]
  assign HanningBlock_io_HanningSignal_ready = FFTBlock_io_din_ready; // @[STFT.scala 35:39]
  assign FFTBlock_clock = clock;
  assign FFTBlock_reset = reset;
  assign FFTBlock_io_din_valid = HanningBlock_io_HanningSignal_valid; // @[STFT.scala 34:25]
  assign FFTBlock_io_din_bits_re = HanningBlock_io_HanningSignal_bits_value; // @[STFT.scala 33:24]
  assign FFTBlock_io_dout_ready = SpectrogramGenBlock_io_FFTsignal_ready; // @[STFT.scala 37:20]
  assign SpectrogramGenBlock_clock = clock;
  assign SpectrogramGenBlock_reset = reset;
  assign SpectrogramGenBlock_io_FFTsignal_valid = FFTBlock_io_dout_valid; // @[STFT.scala 37:20]
  assign SpectrogramGenBlock_io_FFTsignal_bits_re = FFTBlock_io_dout_bits_re; // @[STFT.scala 37:20]
  assign SpectrogramGenBlock_io_FFTsignal_bits_im = FFTBlock_io_dout_bits_im; // @[STFT.scala 37:20]
  assign SpectrogramGenBlock_io_Spectrogram_ready = io_spectrogram_ready; // @[STFT.scala 39:18]
endmodule
