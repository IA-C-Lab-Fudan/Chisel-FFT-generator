module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T; // @[Butterfly.scala 57:28]
  wire [63:0] _T_1; // @[Butterfly.scala 57:52]
  wire [63:0] _T_4; // @[Butterfly.scala 57:40]
  wire [63:0] _T_5; // @[Butterfly.scala 58:28]
  wire [63:0] _T_6; // @[Butterfly.scala 58:52]
  wire [63:0] _T_9; // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2; // @[Butterfly.scala 58:15]
  assign _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  assign _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  assign _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  assign _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  assign _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  assign _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  assign _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT512(
      input clk_in1_p,
    input clk_in1_n,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
    wire clock;
    clk_wiz_0 clk_wiz_0_inst0
       (
        // Clock out ports
        .clk_out1(clock),     // output clk_out1
       // Clock in ports
        .clk_in1_p(clk_in1_p),    // input clk_in1_p
        .clk_in1_n(clk_in1_n));    // input clk_in1_n
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [8:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [8:0] _T_1; // @[FFT.scala 42:16]
  wire [31:0] _GEN_2; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6; // @[FFT.scala 34:12]
  wire [31:0] _GEN_7; // @[FFT.scala 34:12]
  wire [31:0] _GEN_8; // @[FFT.scala 34:12]
  wire [31:0] _GEN_9; // @[FFT.scala 34:12]
  wire [31:0] _GEN_10; // @[FFT.scala 34:12]
  wire [31:0] _GEN_11; // @[FFT.scala 34:12]
  wire [31:0] _GEN_12; // @[FFT.scala 34:12]
  wire [31:0] _GEN_13; // @[FFT.scala 34:12]
  wire [31:0] _GEN_14; // @[FFT.scala 34:12]
  wire [31:0] _GEN_15; // @[FFT.scala 34:12]
  wire [31:0] _GEN_16; // @[FFT.scala 34:12]
  wire [31:0] _GEN_17; // @[FFT.scala 34:12]
  wire [31:0] _GEN_18; // @[FFT.scala 34:12]
  wire [31:0] _GEN_19; // @[FFT.scala 34:12]
  wire [31:0] _GEN_20; // @[FFT.scala 34:12]
  wire [31:0] _GEN_21; // @[FFT.scala 34:12]
  wire [31:0] _GEN_22; // @[FFT.scala 34:12]
  wire [31:0] _GEN_23; // @[FFT.scala 34:12]
  wire [31:0] _GEN_24; // @[FFT.scala 34:12]
  wire [31:0] _GEN_25; // @[FFT.scala 34:12]
  wire [31:0] _GEN_26; // @[FFT.scala 34:12]
  wire [31:0] _GEN_27; // @[FFT.scala 34:12]
  wire [31:0] _GEN_28; // @[FFT.scala 34:12]
  wire [31:0] _GEN_29; // @[FFT.scala 34:12]
  wire [31:0] _GEN_30; // @[FFT.scala 34:12]
  wire [31:0] _GEN_31; // @[FFT.scala 34:12]
  wire [31:0] _GEN_32; // @[FFT.scala 34:12]
  wire [31:0] _GEN_33; // @[FFT.scala 34:12]
  wire [31:0] _GEN_34; // @[FFT.scala 34:12]
  wire [31:0] _GEN_35; // @[FFT.scala 34:12]
  wire [31:0] _GEN_36; // @[FFT.scala 34:12]
  wire [31:0] _GEN_37; // @[FFT.scala 34:12]
  wire [31:0] _GEN_38; // @[FFT.scala 34:12]
  wire [31:0] _GEN_39; // @[FFT.scala 34:12]
  wire [31:0] _GEN_40; // @[FFT.scala 34:12]
  wire [31:0] _GEN_41; // @[FFT.scala 34:12]
  wire [31:0] _GEN_42; // @[FFT.scala 34:12]
  wire [31:0] _GEN_43; // @[FFT.scala 34:12]
  wire [31:0] _GEN_44; // @[FFT.scala 34:12]
  wire [31:0] _GEN_45; // @[FFT.scala 34:12]
  wire [31:0] _GEN_46; // @[FFT.scala 34:12]
  wire [31:0] _GEN_47; // @[FFT.scala 34:12]
  wire [31:0] _GEN_48; // @[FFT.scala 34:12]
  wire [31:0] _GEN_49; // @[FFT.scala 34:12]
  wire [31:0] _GEN_50; // @[FFT.scala 34:12]
  wire [31:0] _GEN_51; // @[FFT.scala 34:12]
  wire [31:0] _GEN_52; // @[FFT.scala 34:12]
  wire [31:0] _GEN_53; // @[FFT.scala 34:12]
  wire [31:0] _GEN_54; // @[FFT.scala 34:12]
  wire [31:0] _GEN_55; // @[FFT.scala 34:12]
  wire [31:0] _GEN_56; // @[FFT.scala 34:12]
  wire [31:0] _GEN_57; // @[FFT.scala 34:12]
  wire [31:0] _GEN_58; // @[FFT.scala 34:12]
  wire [31:0] _GEN_59; // @[FFT.scala 34:12]
  wire [31:0] _GEN_60; // @[FFT.scala 34:12]
  wire [31:0] _GEN_61; // @[FFT.scala 34:12]
  wire [31:0] _GEN_62; // @[FFT.scala 34:12]
  wire [31:0] _GEN_63; // @[FFT.scala 34:12]
  wire [31:0] _GEN_64; // @[FFT.scala 34:12]
  wire [31:0] _GEN_65; // @[FFT.scala 34:12]
  wire [31:0] _GEN_66; // @[FFT.scala 34:12]
  wire [31:0] _GEN_67; // @[FFT.scala 34:12]
  wire [31:0] _GEN_68; // @[FFT.scala 34:12]
  wire [31:0] _GEN_69; // @[FFT.scala 34:12]
  wire [31:0] _GEN_70; // @[FFT.scala 34:12]
  wire [31:0] _GEN_71; // @[FFT.scala 34:12]
  wire [31:0] _GEN_72; // @[FFT.scala 34:12]
  wire [31:0] _GEN_73; // @[FFT.scala 34:12]
  wire [31:0] _GEN_74; // @[FFT.scala 34:12]
  wire [31:0] _GEN_75; // @[FFT.scala 34:12]
  wire [31:0] _GEN_76; // @[FFT.scala 34:12]
  wire [31:0] _GEN_77; // @[FFT.scala 34:12]
  wire [31:0] _GEN_78; // @[FFT.scala 34:12]
  wire [31:0] _GEN_79; // @[FFT.scala 34:12]
  wire [31:0] _GEN_80; // @[FFT.scala 34:12]
  wire [31:0] _GEN_81; // @[FFT.scala 34:12]
  wire [31:0] _GEN_82; // @[FFT.scala 34:12]
  wire [31:0] _GEN_83; // @[FFT.scala 34:12]
  wire [31:0] _GEN_84; // @[FFT.scala 34:12]
  wire [31:0] _GEN_85; // @[FFT.scala 34:12]
  wire [31:0] _GEN_86; // @[FFT.scala 34:12]
  wire [31:0] _GEN_87; // @[FFT.scala 34:12]
  wire [31:0] _GEN_88; // @[FFT.scala 34:12]
  wire [31:0] _GEN_89; // @[FFT.scala 34:12]
  wire [31:0] _GEN_90; // @[FFT.scala 34:12]
  wire [31:0] _GEN_91; // @[FFT.scala 34:12]
  wire [31:0] _GEN_92; // @[FFT.scala 34:12]
  wire [31:0] _GEN_93; // @[FFT.scala 34:12]
  wire [31:0] _GEN_94; // @[FFT.scala 34:12]
  wire [31:0] _GEN_95; // @[FFT.scala 34:12]
  wire [31:0] _GEN_96; // @[FFT.scala 34:12]
  wire [31:0] _GEN_97; // @[FFT.scala 34:12]
  wire [31:0] _GEN_98; // @[FFT.scala 34:12]
  wire [31:0] _GEN_99; // @[FFT.scala 34:12]
  wire [31:0] _GEN_100; // @[FFT.scala 34:12]
  wire [31:0] _GEN_101; // @[FFT.scala 34:12]
  wire [31:0] _GEN_102; // @[FFT.scala 34:12]
  wire [31:0] _GEN_103; // @[FFT.scala 34:12]
  wire [31:0] _GEN_104; // @[FFT.scala 34:12]
  wire [31:0] _GEN_105; // @[FFT.scala 34:12]
  wire [31:0] _GEN_106; // @[FFT.scala 34:12]
  wire [31:0] _GEN_107; // @[FFT.scala 34:12]
  wire [31:0] _GEN_108; // @[FFT.scala 34:12]
  wire [31:0] _GEN_109; // @[FFT.scala 34:12]
  wire [31:0] _GEN_110; // @[FFT.scala 34:12]
  wire [31:0] _GEN_111; // @[FFT.scala 34:12]
  wire [31:0] _GEN_112; // @[FFT.scala 34:12]
  wire [31:0] _GEN_113; // @[FFT.scala 34:12]
  wire [31:0] _GEN_114; // @[FFT.scala 34:12]
  wire [31:0] _GEN_115; // @[FFT.scala 34:12]
  wire [31:0] _GEN_116; // @[FFT.scala 34:12]
  wire [31:0] _GEN_117; // @[FFT.scala 34:12]
  wire [31:0] _GEN_118; // @[FFT.scala 34:12]
  wire [31:0] _GEN_119; // @[FFT.scala 34:12]
  wire [31:0] _GEN_120; // @[FFT.scala 34:12]
  wire [31:0] _GEN_121; // @[FFT.scala 34:12]
  wire [31:0] _GEN_122; // @[FFT.scala 34:12]
  wire [31:0] _GEN_123; // @[FFT.scala 34:12]
  wire [31:0] _GEN_124; // @[FFT.scala 34:12]
  wire [31:0] _GEN_125; // @[FFT.scala 34:12]
  wire [31:0] _GEN_126; // @[FFT.scala 34:12]
  wire [31:0] _GEN_127; // @[FFT.scala 34:12]
  wire [31:0] _GEN_128; // @[FFT.scala 34:12]
  wire [31:0] _GEN_129; // @[FFT.scala 34:12]
  wire [31:0] _GEN_130; // @[FFT.scala 34:12]
  wire [31:0] _GEN_131; // @[FFT.scala 34:12]
  wire [31:0] _GEN_132; // @[FFT.scala 34:12]
  wire [31:0] _GEN_133; // @[FFT.scala 34:12]
  wire [31:0] _GEN_134; // @[FFT.scala 34:12]
  wire [31:0] _GEN_135; // @[FFT.scala 34:12]
  wire [31:0] _GEN_136; // @[FFT.scala 34:12]
  wire [31:0] _GEN_137; // @[FFT.scala 34:12]
  wire [31:0] _GEN_138; // @[FFT.scala 34:12]
  wire [31:0] _GEN_139; // @[FFT.scala 34:12]
  wire [31:0] _GEN_140; // @[FFT.scala 34:12]
  wire [31:0] _GEN_141; // @[FFT.scala 34:12]
  wire [31:0] _GEN_142; // @[FFT.scala 34:12]
  wire [31:0] _GEN_143; // @[FFT.scala 34:12]
  wire [31:0] _GEN_144; // @[FFT.scala 34:12]
  wire [31:0] _GEN_145; // @[FFT.scala 34:12]
  wire [31:0] _GEN_146; // @[FFT.scala 34:12]
  wire [31:0] _GEN_147; // @[FFT.scala 34:12]
  wire [31:0] _GEN_148; // @[FFT.scala 34:12]
  wire [31:0] _GEN_149; // @[FFT.scala 34:12]
  wire [31:0] _GEN_150; // @[FFT.scala 34:12]
  wire [31:0] _GEN_151; // @[FFT.scala 34:12]
  wire [31:0] _GEN_152; // @[FFT.scala 34:12]
  wire [31:0] _GEN_153; // @[FFT.scala 34:12]
  wire [31:0] _GEN_154; // @[FFT.scala 34:12]
  wire [31:0] _GEN_155; // @[FFT.scala 34:12]
  wire [31:0] _GEN_156; // @[FFT.scala 34:12]
  wire [31:0] _GEN_157; // @[FFT.scala 34:12]
  wire [31:0] _GEN_158; // @[FFT.scala 34:12]
  wire [31:0] _GEN_159; // @[FFT.scala 34:12]
  wire [31:0] _GEN_160; // @[FFT.scala 34:12]
  wire [31:0] _GEN_161; // @[FFT.scala 34:12]
  wire [31:0] _GEN_162; // @[FFT.scala 34:12]
  wire [31:0] _GEN_163; // @[FFT.scala 34:12]
  wire [31:0] _GEN_164; // @[FFT.scala 34:12]
  wire [31:0] _GEN_165; // @[FFT.scala 34:12]
  wire [31:0] _GEN_166; // @[FFT.scala 34:12]
  wire [31:0] _GEN_167; // @[FFT.scala 34:12]
  wire [31:0] _GEN_168; // @[FFT.scala 34:12]
  wire [31:0] _GEN_169; // @[FFT.scala 34:12]
  wire [31:0] _GEN_170; // @[FFT.scala 34:12]
  wire [31:0] _GEN_171; // @[FFT.scala 34:12]
  wire [31:0] _GEN_172; // @[FFT.scala 34:12]
  wire [31:0] _GEN_173; // @[FFT.scala 34:12]
  wire [31:0] _GEN_174; // @[FFT.scala 34:12]
  wire [31:0] _GEN_175; // @[FFT.scala 34:12]
  wire [31:0] _GEN_176; // @[FFT.scala 34:12]
  wire [31:0] _GEN_177; // @[FFT.scala 34:12]
  wire [31:0] _GEN_178; // @[FFT.scala 34:12]
  wire [31:0] _GEN_179; // @[FFT.scala 34:12]
  wire [31:0] _GEN_180; // @[FFT.scala 34:12]
  wire [31:0] _GEN_181; // @[FFT.scala 34:12]
  wire [31:0] _GEN_182; // @[FFT.scala 34:12]
  wire [31:0] _GEN_183; // @[FFT.scala 34:12]
  wire [31:0] _GEN_184; // @[FFT.scala 34:12]
  wire [31:0] _GEN_185; // @[FFT.scala 34:12]
  wire [31:0] _GEN_186; // @[FFT.scala 34:12]
  wire [31:0] _GEN_187; // @[FFT.scala 34:12]
  wire [31:0] _GEN_188; // @[FFT.scala 34:12]
  wire [31:0] _GEN_189; // @[FFT.scala 34:12]
  wire [31:0] _GEN_190; // @[FFT.scala 34:12]
  wire [31:0] _GEN_191; // @[FFT.scala 34:12]
  wire [31:0] _GEN_192; // @[FFT.scala 34:12]
  wire [31:0] _GEN_193; // @[FFT.scala 34:12]
  wire [31:0] _GEN_194; // @[FFT.scala 34:12]
  wire [31:0] _GEN_195; // @[FFT.scala 34:12]
  wire [31:0] _GEN_196; // @[FFT.scala 34:12]
  wire [31:0] _GEN_197; // @[FFT.scala 34:12]
  wire [31:0] _GEN_198; // @[FFT.scala 34:12]
  wire [31:0] _GEN_199; // @[FFT.scala 34:12]
  wire [31:0] _GEN_200; // @[FFT.scala 34:12]
  wire [31:0] _GEN_201; // @[FFT.scala 34:12]
  wire [31:0] _GEN_202; // @[FFT.scala 34:12]
  wire [31:0] _GEN_203; // @[FFT.scala 34:12]
  wire [31:0] _GEN_204; // @[FFT.scala 34:12]
  wire [31:0] _GEN_205; // @[FFT.scala 34:12]
  wire [31:0] _GEN_206; // @[FFT.scala 34:12]
  wire [31:0] _GEN_207; // @[FFT.scala 34:12]
  wire [31:0] _GEN_208; // @[FFT.scala 34:12]
  wire [31:0] _GEN_209; // @[FFT.scala 34:12]
  wire [31:0] _GEN_210; // @[FFT.scala 34:12]
  wire [31:0] _GEN_211; // @[FFT.scala 34:12]
  wire [31:0] _GEN_212; // @[FFT.scala 34:12]
  wire [31:0] _GEN_213; // @[FFT.scala 34:12]
  wire [31:0] _GEN_214; // @[FFT.scala 34:12]
  wire [31:0] _GEN_215; // @[FFT.scala 34:12]
  wire [31:0] _GEN_216; // @[FFT.scala 34:12]
  wire [31:0] _GEN_217; // @[FFT.scala 34:12]
  wire [31:0] _GEN_218; // @[FFT.scala 34:12]
  wire [31:0] _GEN_219; // @[FFT.scala 34:12]
  wire [31:0] _GEN_220; // @[FFT.scala 34:12]
  wire [31:0] _GEN_221; // @[FFT.scala 34:12]
  wire [31:0] _GEN_222; // @[FFT.scala 34:12]
  wire [31:0] _GEN_223; // @[FFT.scala 34:12]
  wire [31:0] _GEN_224; // @[FFT.scala 34:12]
  wire [31:0] _GEN_225; // @[FFT.scala 34:12]
  wire [31:0] _GEN_226; // @[FFT.scala 34:12]
  wire [31:0] _GEN_227; // @[FFT.scala 34:12]
  wire [31:0] _GEN_228; // @[FFT.scala 34:12]
  wire [31:0] _GEN_229; // @[FFT.scala 34:12]
  wire [31:0] _GEN_230; // @[FFT.scala 34:12]
  wire [31:0] _GEN_231; // @[FFT.scala 34:12]
  wire [31:0] _GEN_232; // @[FFT.scala 34:12]
  wire [31:0] _GEN_233; // @[FFT.scala 34:12]
  wire [31:0] _GEN_234; // @[FFT.scala 34:12]
  wire [31:0] _GEN_235; // @[FFT.scala 34:12]
  wire [31:0] _GEN_236; // @[FFT.scala 34:12]
  wire [31:0] _GEN_237; // @[FFT.scala 34:12]
  wire [31:0] _GEN_238; // @[FFT.scala 34:12]
  wire [31:0] _GEN_239; // @[FFT.scala 34:12]
  wire [31:0] _GEN_240; // @[FFT.scala 34:12]
  wire [31:0] _GEN_241; // @[FFT.scala 34:12]
  wire [31:0] _GEN_242; // @[FFT.scala 34:12]
  wire [31:0] _GEN_243; // @[FFT.scala 34:12]
  wire [31:0] _GEN_244; // @[FFT.scala 34:12]
  wire [31:0] _GEN_245; // @[FFT.scala 34:12]
  wire [31:0] _GEN_246; // @[FFT.scala 34:12]
  wire [31:0] _GEN_247; // @[FFT.scala 34:12]
  wire [31:0] _GEN_248; // @[FFT.scala 34:12]
  wire [31:0] _GEN_249; // @[FFT.scala 34:12]
  wire [31:0] _GEN_250; // @[FFT.scala 34:12]
  wire [31:0] _GEN_251; // @[FFT.scala 34:12]
  wire [31:0] _GEN_252; // @[FFT.scala 34:12]
  wire [31:0] _GEN_253; // @[FFT.scala 34:12]
  wire [31:0] _GEN_254; // @[FFT.scala 34:12]
  wire [31:0] _GEN_255; // @[FFT.scala 34:12]
  wire [31:0] _GEN_258; // @[FFT.scala 35:12]
  wire [31:0] _GEN_259; // @[FFT.scala 35:12]
  wire [31:0] _GEN_260; // @[FFT.scala 35:12]
  wire [31:0] _GEN_261; // @[FFT.scala 35:12]
  wire [31:0] _GEN_262; // @[FFT.scala 35:12]
  wire [31:0] _GEN_263; // @[FFT.scala 35:12]
  wire [31:0] _GEN_264; // @[FFT.scala 35:12]
  wire [31:0] _GEN_265; // @[FFT.scala 35:12]
  wire [31:0] _GEN_266; // @[FFT.scala 35:12]
  wire [31:0] _GEN_267; // @[FFT.scala 35:12]
  wire [31:0] _GEN_268; // @[FFT.scala 35:12]
  wire [31:0] _GEN_269; // @[FFT.scala 35:12]
  wire [31:0] _GEN_270; // @[FFT.scala 35:12]
  wire [31:0] _GEN_271; // @[FFT.scala 35:12]
  wire [31:0] _GEN_272; // @[FFT.scala 35:12]
  wire [31:0] _GEN_273; // @[FFT.scala 35:12]
  wire [31:0] _GEN_274; // @[FFT.scala 35:12]
  wire [31:0] _GEN_275; // @[FFT.scala 35:12]
  wire [31:0] _GEN_276; // @[FFT.scala 35:12]
  wire [31:0] _GEN_277; // @[FFT.scala 35:12]
  wire [31:0] _GEN_278; // @[FFT.scala 35:12]
  wire [31:0] _GEN_279; // @[FFT.scala 35:12]
  wire [31:0] _GEN_280; // @[FFT.scala 35:12]
  wire [31:0] _GEN_281; // @[FFT.scala 35:12]
  wire [31:0] _GEN_282; // @[FFT.scala 35:12]
  wire [31:0] _GEN_283; // @[FFT.scala 35:12]
  wire [31:0] _GEN_284; // @[FFT.scala 35:12]
  wire [31:0] _GEN_285; // @[FFT.scala 35:12]
  wire [31:0] _GEN_286; // @[FFT.scala 35:12]
  wire [31:0] _GEN_287; // @[FFT.scala 35:12]
  wire [31:0] _GEN_288; // @[FFT.scala 35:12]
  wire [31:0] _GEN_289; // @[FFT.scala 35:12]
  wire [31:0] _GEN_290; // @[FFT.scala 35:12]
  wire [31:0] _GEN_291; // @[FFT.scala 35:12]
  wire [31:0] _GEN_292; // @[FFT.scala 35:12]
  wire [31:0] _GEN_293; // @[FFT.scala 35:12]
  wire [31:0] _GEN_294; // @[FFT.scala 35:12]
  wire [31:0] _GEN_295; // @[FFT.scala 35:12]
  wire [31:0] _GEN_296; // @[FFT.scala 35:12]
  wire [31:0] _GEN_297; // @[FFT.scala 35:12]
  wire [31:0] _GEN_298; // @[FFT.scala 35:12]
  wire [31:0] _GEN_299; // @[FFT.scala 35:12]
  wire [31:0] _GEN_300; // @[FFT.scala 35:12]
  wire [31:0] _GEN_301; // @[FFT.scala 35:12]
  wire [31:0] _GEN_302; // @[FFT.scala 35:12]
  wire [31:0] _GEN_303; // @[FFT.scala 35:12]
  wire [31:0] _GEN_304; // @[FFT.scala 35:12]
  wire [31:0] _GEN_305; // @[FFT.scala 35:12]
  wire [31:0] _GEN_306; // @[FFT.scala 35:12]
  wire [31:0] _GEN_307; // @[FFT.scala 35:12]
  wire [31:0] _GEN_308; // @[FFT.scala 35:12]
  wire [31:0] _GEN_309; // @[FFT.scala 35:12]
  wire [31:0] _GEN_310; // @[FFT.scala 35:12]
  wire [31:0] _GEN_311; // @[FFT.scala 35:12]
  wire [31:0] _GEN_312; // @[FFT.scala 35:12]
  wire [31:0] _GEN_313; // @[FFT.scala 35:12]
  wire [31:0] _GEN_314; // @[FFT.scala 35:12]
  wire [31:0] _GEN_315; // @[FFT.scala 35:12]
  wire [31:0] _GEN_316; // @[FFT.scala 35:12]
  wire [31:0] _GEN_317; // @[FFT.scala 35:12]
  wire [31:0] _GEN_318; // @[FFT.scala 35:12]
  wire [31:0] _GEN_319; // @[FFT.scala 35:12]
  wire [31:0] _GEN_320; // @[FFT.scala 35:12]
  wire [31:0] _GEN_321; // @[FFT.scala 35:12]
  wire [31:0] _GEN_322; // @[FFT.scala 35:12]
  wire [31:0] _GEN_323; // @[FFT.scala 35:12]
  wire [31:0] _GEN_324; // @[FFT.scala 35:12]
  wire [31:0] _GEN_325; // @[FFT.scala 35:12]
  wire [31:0] _GEN_326; // @[FFT.scala 35:12]
  wire [31:0] _GEN_327; // @[FFT.scala 35:12]
  wire [31:0] _GEN_328; // @[FFT.scala 35:12]
  wire [31:0] _GEN_329; // @[FFT.scala 35:12]
  wire [31:0] _GEN_330; // @[FFT.scala 35:12]
  wire [31:0] _GEN_331; // @[FFT.scala 35:12]
  wire [31:0] _GEN_332; // @[FFT.scala 35:12]
  wire [31:0] _GEN_333; // @[FFT.scala 35:12]
  wire [31:0] _GEN_334; // @[FFT.scala 35:12]
  wire [31:0] _GEN_335; // @[FFT.scala 35:12]
  wire [31:0] _GEN_336; // @[FFT.scala 35:12]
  wire [31:0] _GEN_337; // @[FFT.scala 35:12]
  wire [31:0] _GEN_338; // @[FFT.scala 35:12]
  wire [31:0] _GEN_339; // @[FFT.scala 35:12]
  wire [31:0] _GEN_340; // @[FFT.scala 35:12]
  wire [31:0] _GEN_341; // @[FFT.scala 35:12]
  wire [31:0] _GEN_342; // @[FFT.scala 35:12]
  wire [31:0] _GEN_343; // @[FFT.scala 35:12]
  wire [31:0] _GEN_344; // @[FFT.scala 35:12]
  wire [31:0] _GEN_345; // @[FFT.scala 35:12]
  wire [31:0] _GEN_346; // @[FFT.scala 35:12]
  wire [31:0] _GEN_347; // @[FFT.scala 35:12]
  wire [31:0] _GEN_348; // @[FFT.scala 35:12]
  wire [31:0] _GEN_349; // @[FFT.scala 35:12]
  wire [31:0] _GEN_350; // @[FFT.scala 35:12]
  wire [31:0] _GEN_351; // @[FFT.scala 35:12]
  wire [31:0] _GEN_352; // @[FFT.scala 35:12]
  wire [31:0] _GEN_353; // @[FFT.scala 35:12]
  wire [31:0] _GEN_354; // @[FFT.scala 35:12]
  wire [31:0] _GEN_355; // @[FFT.scala 35:12]
  wire [31:0] _GEN_356; // @[FFT.scala 35:12]
  wire [31:0] _GEN_357; // @[FFT.scala 35:12]
  wire [31:0] _GEN_358; // @[FFT.scala 35:12]
  wire [31:0] _GEN_359; // @[FFT.scala 35:12]
  wire [31:0] _GEN_360; // @[FFT.scala 35:12]
  wire [31:0] _GEN_361; // @[FFT.scala 35:12]
  wire [31:0] _GEN_362; // @[FFT.scala 35:12]
  wire [31:0] _GEN_363; // @[FFT.scala 35:12]
  wire [31:0] _GEN_364; // @[FFT.scala 35:12]
  wire [31:0] _GEN_365; // @[FFT.scala 35:12]
  wire [31:0] _GEN_366; // @[FFT.scala 35:12]
  wire [31:0] _GEN_367; // @[FFT.scala 35:12]
  wire [31:0] _GEN_368; // @[FFT.scala 35:12]
  wire [31:0] _GEN_369; // @[FFT.scala 35:12]
  wire [31:0] _GEN_370; // @[FFT.scala 35:12]
  wire [31:0] _GEN_371; // @[FFT.scala 35:12]
  wire [31:0] _GEN_372; // @[FFT.scala 35:12]
  wire [31:0] _GEN_373; // @[FFT.scala 35:12]
  wire [31:0] _GEN_374; // @[FFT.scala 35:12]
  wire [31:0] _GEN_375; // @[FFT.scala 35:12]
  wire [31:0] _GEN_376; // @[FFT.scala 35:12]
  wire [31:0] _GEN_377; // @[FFT.scala 35:12]
  wire [31:0] _GEN_378; // @[FFT.scala 35:12]
  wire [31:0] _GEN_379; // @[FFT.scala 35:12]
  wire [31:0] _GEN_380; // @[FFT.scala 35:12]
  wire [31:0] _GEN_381; // @[FFT.scala 35:12]
  wire [31:0] _GEN_382; // @[FFT.scala 35:12]
  wire [31:0] _GEN_383; // @[FFT.scala 35:12]
  wire [31:0] _GEN_384; // @[FFT.scala 35:12]
  wire [31:0] _GEN_385; // @[FFT.scala 35:12]
  wire [31:0] _GEN_386; // @[FFT.scala 35:12]
  wire [31:0] _GEN_387; // @[FFT.scala 35:12]
  wire [31:0] _GEN_388; // @[FFT.scala 35:12]
  wire [31:0] _GEN_389; // @[FFT.scala 35:12]
  wire [31:0] _GEN_390; // @[FFT.scala 35:12]
  wire [31:0] _GEN_391; // @[FFT.scala 35:12]
  wire [31:0] _GEN_392; // @[FFT.scala 35:12]
  wire [31:0] _GEN_393; // @[FFT.scala 35:12]
  wire [31:0] _GEN_394; // @[FFT.scala 35:12]
  wire [31:0] _GEN_395; // @[FFT.scala 35:12]
  wire [31:0] _GEN_396; // @[FFT.scala 35:12]
  wire [31:0] _GEN_397; // @[FFT.scala 35:12]
  wire [31:0] _GEN_398; // @[FFT.scala 35:12]
  wire [31:0] _GEN_399; // @[FFT.scala 35:12]
  wire [31:0] _GEN_400; // @[FFT.scala 35:12]
  wire [31:0] _GEN_401; // @[FFT.scala 35:12]
  wire [31:0] _GEN_402; // @[FFT.scala 35:12]
  wire [31:0] _GEN_403; // @[FFT.scala 35:12]
  wire [31:0] _GEN_404; // @[FFT.scala 35:12]
  wire [31:0] _GEN_405; // @[FFT.scala 35:12]
  wire [31:0] _GEN_406; // @[FFT.scala 35:12]
  wire [31:0] _GEN_407; // @[FFT.scala 35:12]
  wire [31:0] _GEN_408; // @[FFT.scala 35:12]
  wire [31:0] _GEN_409; // @[FFT.scala 35:12]
  wire [31:0] _GEN_410; // @[FFT.scala 35:12]
  wire [31:0] _GEN_411; // @[FFT.scala 35:12]
  wire [31:0] _GEN_412; // @[FFT.scala 35:12]
  wire [31:0] _GEN_413; // @[FFT.scala 35:12]
  wire [31:0] _GEN_414; // @[FFT.scala 35:12]
  wire [31:0] _GEN_415; // @[FFT.scala 35:12]
  wire [31:0] _GEN_416; // @[FFT.scala 35:12]
  wire [31:0] _GEN_417; // @[FFT.scala 35:12]
  wire [31:0] _GEN_418; // @[FFT.scala 35:12]
  wire [31:0] _GEN_419; // @[FFT.scala 35:12]
  wire [31:0] _GEN_420; // @[FFT.scala 35:12]
  wire [31:0] _GEN_421; // @[FFT.scala 35:12]
  wire [31:0] _GEN_422; // @[FFT.scala 35:12]
  wire [31:0] _GEN_423; // @[FFT.scala 35:12]
  wire [31:0] _GEN_424; // @[FFT.scala 35:12]
  wire [31:0] _GEN_425; // @[FFT.scala 35:12]
  wire [31:0] _GEN_426; // @[FFT.scala 35:12]
  wire [31:0] _GEN_427; // @[FFT.scala 35:12]
  wire [31:0] _GEN_428; // @[FFT.scala 35:12]
  wire [31:0] _GEN_429; // @[FFT.scala 35:12]
  wire [31:0] _GEN_430; // @[FFT.scala 35:12]
  wire [31:0] _GEN_431; // @[FFT.scala 35:12]
  wire [31:0] _GEN_432; // @[FFT.scala 35:12]
  wire [31:0] _GEN_433; // @[FFT.scala 35:12]
  wire [31:0] _GEN_434; // @[FFT.scala 35:12]
  wire [31:0] _GEN_435; // @[FFT.scala 35:12]
  wire [31:0] _GEN_436; // @[FFT.scala 35:12]
  wire [31:0] _GEN_437; // @[FFT.scala 35:12]
  wire [31:0] _GEN_438; // @[FFT.scala 35:12]
  wire [31:0] _GEN_439; // @[FFT.scala 35:12]
  wire [31:0] _GEN_440; // @[FFT.scala 35:12]
  wire [31:0] _GEN_441; // @[FFT.scala 35:12]
  wire [31:0] _GEN_442; // @[FFT.scala 35:12]
  wire [31:0] _GEN_443; // @[FFT.scala 35:12]
  wire [31:0] _GEN_444; // @[FFT.scala 35:12]
  wire [31:0] _GEN_445; // @[FFT.scala 35:12]
  wire [31:0] _GEN_446; // @[FFT.scala 35:12]
  wire [31:0] _GEN_447; // @[FFT.scala 35:12]
  wire [31:0] _GEN_448; // @[FFT.scala 35:12]
  wire [31:0] _GEN_449; // @[FFT.scala 35:12]
  wire [31:0] _GEN_450; // @[FFT.scala 35:12]
  wire [31:0] _GEN_451; // @[FFT.scala 35:12]
  wire [31:0] _GEN_452; // @[FFT.scala 35:12]
  wire [31:0] _GEN_453; // @[FFT.scala 35:12]
  wire [31:0] _GEN_454; // @[FFT.scala 35:12]
  wire [31:0] _GEN_455; // @[FFT.scala 35:12]
  wire [31:0] _GEN_456; // @[FFT.scala 35:12]
  wire [31:0] _GEN_457; // @[FFT.scala 35:12]
  wire [31:0] _GEN_458; // @[FFT.scala 35:12]
  wire [31:0] _GEN_459; // @[FFT.scala 35:12]
  wire [31:0] _GEN_460; // @[FFT.scala 35:12]
  wire [31:0] _GEN_461; // @[FFT.scala 35:12]
  wire [31:0] _GEN_462; // @[FFT.scala 35:12]
  wire [31:0] _GEN_463; // @[FFT.scala 35:12]
  wire [31:0] _GEN_464; // @[FFT.scala 35:12]
  wire [31:0] _GEN_465; // @[FFT.scala 35:12]
  wire [31:0] _GEN_466; // @[FFT.scala 35:12]
  wire [31:0] _GEN_467; // @[FFT.scala 35:12]
  wire [31:0] _GEN_468; // @[FFT.scala 35:12]
  wire [31:0] _GEN_469; // @[FFT.scala 35:12]
  wire [31:0] _GEN_470; // @[FFT.scala 35:12]
  wire [31:0] _GEN_471; // @[FFT.scala 35:12]
  wire [31:0] _GEN_472; // @[FFT.scala 35:12]
  wire [31:0] _GEN_473; // @[FFT.scala 35:12]
  wire [31:0] _GEN_474; // @[FFT.scala 35:12]
  wire [31:0] _GEN_475; // @[FFT.scala 35:12]
  wire [31:0] _GEN_476; // @[FFT.scala 35:12]
  wire [31:0] _GEN_477; // @[FFT.scala 35:12]
  wire [31:0] _GEN_478; // @[FFT.scala 35:12]
  wire [31:0] _GEN_479; // @[FFT.scala 35:12]
  wire [31:0] _GEN_480; // @[FFT.scala 35:12]
  wire [31:0] _GEN_481; // @[FFT.scala 35:12]
  wire [31:0] _GEN_482; // @[FFT.scala 35:12]
  wire [31:0] _GEN_483; // @[FFT.scala 35:12]
  wire [31:0] _GEN_484; // @[FFT.scala 35:12]
  wire [31:0] _GEN_485; // @[FFT.scala 35:12]
  wire [31:0] _GEN_486; // @[FFT.scala 35:12]
  wire [31:0] _GEN_487; // @[FFT.scala 35:12]
  wire [31:0] _GEN_488; // @[FFT.scala 35:12]
  wire [31:0] _GEN_489; // @[FFT.scala 35:12]
  wire [31:0] _GEN_490; // @[FFT.scala 35:12]
  wire [31:0] _GEN_491; // @[FFT.scala 35:12]
  wire [31:0] _GEN_492; // @[FFT.scala 35:12]
  wire [31:0] _GEN_493; // @[FFT.scala 35:12]
  wire [31:0] _GEN_494; // @[FFT.scala 35:12]
  wire [31:0] _GEN_495; // @[FFT.scala 35:12]
  wire [31:0] _GEN_496; // @[FFT.scala 35:12]
  wire [31:0] _GEN_497; // @[FFT.scala 35:12]
  wire [31:0] _GEN_498; // @[FFT.scala 35:12]
  wire [31:0] _GEN_499; // @[FFT.scala 35:12]
  wire [31:0] _GEN_500; // @[FFT.scala 35:12]
  wire [31:0] _GEN_501; // @[FFT.scala 35:12]
  wire [31:0] _GEN_502; // @[FFT.scala 35:12]
  wire [31:0] _GEN_503; // @[FFT.scala 35:12]
  wire [31:0] _GEN_504; // @[FFT.scala 35:12]
  wire [31:0] _GEN_505; // @[FFT.scala 35:12]
  wire [31:0] _GEN_506; // @[FFT.scala 35:12]
  wire [31:0] _GEN_507; // @[FFT.scala 35:12]
  wire [31:0] _GEN_508; // @[FFT.scala 35:12]
  wire [31:0] _GEN_509; // @[FFT.scala 35:12]
  wire [31:0] _GEN_510; // @[FFT.scala 35:12]
  wire [31:0] _GEN_511; // @[FFT.scala 35:12]
  reg [31:0] _T_146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [31:0] _T_146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [31:0] _T_147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [31:0] _T_147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [31:0] _T_148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [31:0] _T_149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [31:0] _T_393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [31:0] _T_406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_521;
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_522;
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_523;
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_524;
  reg [31:0] _T_409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_525;
  reg [31:0] _T_409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_526;
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_527;
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_528;
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_529;
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_530;
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_531;
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_532;
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_533;
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_534;
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_535;
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_536;
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_537;
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_538;
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_539;
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_540;
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_541;
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_552;
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_553;
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_554;
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_557;
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_558;
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_559;
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_560;
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_561;
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_562;
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_563;
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_564;
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_565;
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_566;
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_567;
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_568;
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_569;
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_570;
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_571;
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_572;
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_573;
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_574;
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_575;
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_576;
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_577;
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_578;
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_579;
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_580;
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_581;
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_582;
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_583;
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_584;
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_585;
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_586;
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_587;
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_588;
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_589;
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_590;
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_591;
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_592;
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_593;
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_594;
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_595;
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_596;
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_597;
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_598;
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_599;
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_600;
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_601;
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_602;
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_603;
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_604;
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_605;
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_606;
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_607;
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_608;
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_609;
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_610;
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_611;
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_612;
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_613;
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_614;
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_615;
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_616;
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_617;
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_618;
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_619;
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_620;
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_621;
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_622;
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_623;
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_624;
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_625;
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_626;
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_627;
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_628;
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_629;
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_630;
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_631;
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_632;
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_633;
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_634;
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_635;
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_636;
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_637;
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_638;
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_639;
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_640;
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_641;
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_642;
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_643;
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_644;
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_645;
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_646;
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_647;
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_648;
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_649;
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_650;
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_651;
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_652;
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_653;
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_654;
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_655;
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_656;
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_657;
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_658;
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_659;
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_660;
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_661;
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_662;
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_663;
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_664;
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_665;
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_666;
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_667;
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_668;
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_669;
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_670;
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_671;
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_672;
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_673;
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_674;
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_675;
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_676;
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_677;
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_678;
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_679;
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_680;
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_681;
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_682;
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_683;
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_684;
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_685;
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_686;
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_687;
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_688;
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_689;
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_690;
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_691;
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_692;
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_693;
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_694;
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_695;
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_696;
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_697;
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_698;
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_699;
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_700;
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_701;
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_702;
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_703;
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_704;
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_705;
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_706;
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_707;
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_708;
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_709;
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_710;
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_711;
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_712;
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_713;
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_714;
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_715;
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_716;
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_717;
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_718;
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_719;
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_720;
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_721;
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_722;
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_723;
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_724;
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_725;
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_726;
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_727;
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_728;
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_729;
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_730;
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_731;
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_732;
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_733;
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_734;
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_735;
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_736;
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_737;
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_738;
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_739;
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_740;
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_741;
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_742;
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_743;
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_744;
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_745;
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_746;
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_747;
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_748;
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_749;
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_750;
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_751;
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_752;
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_753;
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_754;
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_755;
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_756;
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_757;
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_758;
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_759;
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_760;
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_761;
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_762;
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_763;
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_764;
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_765;
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_766;
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_767;
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_768;
  wire [31:0] _GEN_1282; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1283; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1284; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1285; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1286; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1287; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1288; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1289; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1290; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1291; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1292; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1293; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1294; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1295; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1296; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1297; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1298; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1299; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1300; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1301; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1302; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1303; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1304; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1305; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1306; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1307; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1308; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1309; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1310; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1311; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1312; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1313; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1314; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1315; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1316; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1317; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1318; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1319; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1320; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1321; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1322; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1323; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1324; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1325; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1326; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1327; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1328; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1329; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1330; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1331; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1332; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1333; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1334; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1335; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1336; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1337; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1338; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1339; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1340; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1341; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1342; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1343; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1344; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1345; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1346; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1347; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1348; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1349; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1350; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1351; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1352; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1353; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1354; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1355; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1356; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1357; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1358; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1359; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1360; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1361; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1362; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1363; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1364; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1365; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1366; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1367; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1368; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1369; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1370; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1371; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1372; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1373; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1374; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1375; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1376; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1377; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1378; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1379; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1380; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1381; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1382; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1383; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1384; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1385; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1386; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1387; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1388; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1389; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1390; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1391; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1392; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1393; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1394; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1395; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1396; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1397; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1398; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1399; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1400; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1401; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1402; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1403; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1404; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1405; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1406; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1407; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1410; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1411; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1412; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1413; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1414; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1415; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1416; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1417; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1418; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1419; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1420; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1421; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1422; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1423; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1424; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1425; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1426; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1427; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1428; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1429; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1430; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1431; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1432; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1433; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1434; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1435; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1436; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1437; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1438; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1439; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1440; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1441; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1442; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1443; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1444; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1445; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1446; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1447; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1448; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1449; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1450; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1451; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1452; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1453; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1454; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1455; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1456; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1457; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1458; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1459; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1460; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1461; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1462; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1463; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1464; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1465; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1466; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1467; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1468; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1469; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1470; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1471; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1472; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1473; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1474; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1475; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1476; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1477; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1478; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1479; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1480; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1481; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1482; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1483; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1484; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1485; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1486; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1487; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1488; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1489; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1490; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1491; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1492; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1493; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1494; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1495; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1496; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1497; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1498; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1499; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1500; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1501; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1502; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1503; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1504; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1505; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1506; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1507; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1508; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1509; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1510; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1511; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1512; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1513; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1514; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1515; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1516; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1517; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1518; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1519; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1520; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1521; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1522; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1523; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1524; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1525; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1526; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1527; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1528; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1529; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1530; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1531; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1532; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1533; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1534; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1535; // @[FFT.scala 35:12]
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_769;
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  reg [31:0] _T_536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_771;
  reg [31:0] _T_536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_772;
  reg [31:0] _T_537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_773;
  reg [31:0] _T_537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  reg [31:0] _T_538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  reg [31:0] _T_538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  reg [31:0] _T_539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg [31:0] _T_539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  reg [31:0] _T_540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg [31:0] _T_540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  reg [31:0] _T_541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_781;
  reg [31:0] _T_541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_782;
  reg [31:0] _T_542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_783;
  reg [31:0] _T_542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_784;
  reg [31:0] _T_543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_785;
  reg [31:0] _T_543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_786;
  reg [31:0] _T_544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_787;
  reg [31:0] _T_544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_788;
  reg [31:0] _T_545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_789;
  reg [31:0] _T_545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_790;
  reg [31:0] _T_546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_791;
  reg [31:0] _T_546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_792;
  reg [31:0] _T_547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_793;
  reg [31:0] _T_547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_794;
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_795;
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_796;
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_797;
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_798;
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_799;
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_800;
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_801;
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_802;
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_803;
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_804;
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_805;
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_806;
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_807;
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_808;
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_809;
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_810;
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_811;
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_812;
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_813;
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_814;
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_815;
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_816;
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_817;
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_818;
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_819;
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_820;
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_821;
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_822;
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_823;
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_824;
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_825;
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_826;
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_827;
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_828;
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_829;
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_830;
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_831;
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_832;
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_833;
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_834;
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_835;
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_836;
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_837;
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_838;
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_839;
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_840;
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_841;
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_842;
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_843;
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_844;
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_845;
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_846;
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_847;
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_848;
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_849;
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_850;
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_851;
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_852;
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_853;
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_854;
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_855;
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_856;
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_857;
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_858;
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_859;
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_860;
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_861;
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_862;
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_863;
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_864;
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_865;
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_866;
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_867;
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_868;
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_869;
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_870;
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_871;
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_872;
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_873;
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_874;
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_875;
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_876;
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_877;
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_878;
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_879;
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_880;
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_881;
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_882;
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_883;
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_884;
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_885;
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_886;
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_887;
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_888;
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_889;
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_890;
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_891;
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_892;
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_893;
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_894;
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_895;
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_896;
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_897;
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_898;
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_899;
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_900;
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_901;
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_902;
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_903;
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_904;
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_905;
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_906;
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_907;
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_908;
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_909;
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_910;
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_911;
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_912;
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_913;
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_914;
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_915;
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_916;
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_917;
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_918;
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_919;
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_920;
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_921;
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_922;
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_923;
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_924;
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_925;
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_926;
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_927;
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_928;
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_929;
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_930;
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_931;
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_932;
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_933;
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_934;
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_935;
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_936;
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_937;
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_938;
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_939;
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_940;
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_941;
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_942;
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_943;
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_944;
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_945;
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_946;
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_947;
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_948;
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_949;
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_950;
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_951;
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_952;
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_953;
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_954;
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_955;
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_956;
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_957;
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_958;
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_959;
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_960;
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_961;
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_962;
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_963;
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_964;
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_965;
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_966;
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_967;
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_968;
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_969;
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_970;
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_971;
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_972;
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_973;
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_974;
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_975;
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_976;
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_977;
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_978;
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_979;
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_980;
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_981;
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_982;
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_983;
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_984;
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_985;
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_986;
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_987;
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_988;
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_989;
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_990;
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_991;
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_992;
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_993;
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_994;
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_995;
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_996;
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_997;
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_998;
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_999;
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1000;
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1001;
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1002;
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1003;
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1004;
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1005;
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1006;
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1007;
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1008;
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1009;
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1010;
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1011;
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1012;
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1013;
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1014;
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1015;
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1016;
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1017;
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1018;
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1019;
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1020;
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1021;
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1022;
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1023;
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1024;
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1025;
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1026;
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1027;
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1028;
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1029;
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1030;
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1031;
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1032;
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1033;
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1034;
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1035;
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1036;
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1037;
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1038;
  reg [31:0] _T_671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1039;
  reg [31:0] _T_671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1040;
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1041;
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1042;
  reg [31:0] _T_673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1043;
  reg [31:0] _T_673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1044;
  reg [31:0] _T_674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1045;
  reg [31:0] _T_674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1046;
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1047;
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1048;
  reg [31:0] _T_676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1049;
  reg [31:0] _T_676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1050;
  reg [31:0] _T_677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1051;
  reg [31:0] _T_677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1052;
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1053;
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1054;
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1055;
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1056;
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1057;
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1058;
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1059;
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1060;
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1061;
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1062;
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1063;
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1064;
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1065;
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1066;
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1067;
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1068;
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1069;
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1070;
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1071;
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1072;
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1073;
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1074;
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1075;
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1076;
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1077;
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1078;
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1079;
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1080;
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1081;
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1082;
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1083;
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1084;
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1085;
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1086;
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1087;
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1088;
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1089;
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1090;
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1091;
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1092;
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1093;
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1094;
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1095;
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1096;
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1097;
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1098;
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1099;
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1100;
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1101;
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1102;
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1103;
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1104;
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1105;
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1106;
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1107;
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1108;
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1109;
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1110;
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1111;
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1112;
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1113;
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1114;
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1115;
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1116;
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1117;
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1118;
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1119;
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1120;
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1121;
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1122;
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1123;
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1124;
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1125;
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1126;
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1127;
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1128;
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1129;
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1130;
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1131;
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1132;
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1133;
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1134;
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1135;
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1136;
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1137;
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1138;
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1139;
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1140;
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1141;
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1142;
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1143;
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1144;
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1145;
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1146;
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1147;
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1148;
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1149;
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1150;
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1151;
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1152;
  wire [31:0] _GEN_1922; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1923; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1924; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1925; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1926; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1927; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1928; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1929; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1930; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1931; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1932; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1933; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1934; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1935; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1936; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1937; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1938; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1939; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1940; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1941; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1942; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1943; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1944; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1945; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1946; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1947; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1948; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1949; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1950; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1951; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1952; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1953; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1954; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1955; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1956; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1957; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1958; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1959; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1960; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1961; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1962; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1963; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1964; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1965; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1966; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1967; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1968; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1969; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1970; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1971; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1972; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1973; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1974; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1975; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1976; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1977; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1978; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1979; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1980; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1981; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1982; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1983; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1986; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1987; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1988; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1989; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1990; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1991; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1992; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1993; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1994; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1995; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1996; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1997; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1998; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1999; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2000; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2001; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2002; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2003; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2004; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2005; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2006; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2007; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2008; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2009; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2010; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2011; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2012; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2013; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2014; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2015; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2016; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2017; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2018; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2019; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2020; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2021; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2022; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2023; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2024; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2025; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2026; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2027; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2028; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2029; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2030; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2031; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2032; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2033; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2034; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2035; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2036; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2037; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2038; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2039; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2040; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2041; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2042; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2043; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2044; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2045; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2046; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2047; // @[FFT.scala 35:12]
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1153;
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1154;
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1155;
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1156;
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1157;
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1158;
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1159;
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1160;
  reg [31:0] _T_736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1161;
  reg [31:0] _T_736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1162;
  reg [31:0] _T_737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1163;
  reg [31:0] _T_737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1164;
  reg [31:0] _T_738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1165;
  reg [31:0] _T_738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1166;
  reg [31:0] _T_739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1167;
  reg [31:0] _T_739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1168;
  reg [31:0] _T_740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1169;
  reg [31:0] _T_740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1170;
  reg [31:0] _T_741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1171;
  reg [31:0] _T_741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1172;
  reg [31:0] _T_742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1173;
  reg [31:0] _T_742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1174;
  reg [31:0] _T_743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1175;
  reg [31:0] _T_743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1176;
  reg [31:0] _T_744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1177;
  reg [31:0] _T_744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1178;
  reg [31:0] _T_745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1179;
  reg [31:0] _T_745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1180;
  reg [31:0] _T_746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1181;
  reg [31:0] _T_746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1182;
  reg [31:0] _T_747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1183;
  reg [31:0] _T_747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1184;
  reg [31:0] _T_748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1185;
  reg [31:0] _T_748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1186;
  reg [31:0] _T_749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1187;
  reg [31:0] _T_749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1188;
  reg [31:0] _T_750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1189;
  reg [31:0] _T_750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1190;
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1191;
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1192;
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1193;
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1194;
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1195;
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1196;
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1197;
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1198;
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1199;
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1200;
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1201;
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1202;
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1203;
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1204;
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1205;
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1206;
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1207;
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1208;
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1209;
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1210;
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1211;
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1212;
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1213;
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1214;
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1215;
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1216;
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1217;
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1218;
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1219;
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1220;
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1221;
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1222;
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1223;
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1224;
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1225;
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1226;
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1227;
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1228;
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1229;
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1230;
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1231;
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1232;
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1233;
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1234;
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1235;
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1236;
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1237;
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1238;
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1239;
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1240;
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1241;
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1242;
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1243;
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1244;
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1245;
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1246;
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1247;
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1248;
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1249;
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1250;
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1251;
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1252;
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1253;
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1254;
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1255;
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1256;
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1257;
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1258;
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1259;
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1260;
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1261;
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1262;
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1263;
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1264;
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1265;
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1266;
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1267;
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1268;
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1269;
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1270;
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1271;
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1272;
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1273;
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1274;
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1275;
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1276;
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1277;
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1278;
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1279;
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1280;
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1281;
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1282;
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1283;
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1284;
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1285;
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1286;
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1287;
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1288;
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1289;
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1290;
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1291;
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1292;
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1293;
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1294;
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1295;
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1296;
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1297;
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1298;
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1299;
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1300;
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1301;
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1302;
  reg [31:0] _T_808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1303;
  reg [31:0] _T_808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1304;
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1305;
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1306;
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1307;
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1308;
  reg [31:0] _T_811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1309;
  reg [31:0] _T_811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1310;
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1311;
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1312;
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1313;
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1314;
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1315;
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1316;
  reg [31:0] _T_815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1317;
  reg [31:0] _T_815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1318;
  reg [31:0] _T_816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1319;
  reg [31:0] _T_816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1320;
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1321;
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1322;
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1323;
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1324;
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1325;
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1326;
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1327;
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1328;
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1329;
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1330;
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1331;
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1332;
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1333;
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1334;
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1335;
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1336;
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1337;
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1338;
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1339;
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1340;
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1341;
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1342;
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1343;
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1344;
  wire [31:0] _GEN_2242; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2243; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2244; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2245; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2246; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2247; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2248; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2249; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2250; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2251; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2252; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2253; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2254; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2255; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2256; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2257; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2258; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2259; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2260; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2261; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2262; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2263; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2264; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2265; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2266; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2267; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2268; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2269; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2270; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2271; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2274; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2275; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2276; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2277; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2278; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2279; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2280; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2281; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2282; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2283; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2284; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2285; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2286; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2287; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2288; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2289; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2290; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2291; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2292; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2293; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2294; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2295; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2296; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2297; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2298; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2299; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2300; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2301; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2302; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2303; // @[FFT.scala 35:12]
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1345;
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1346;
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1347;
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1348;
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1349;
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1350;
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1351;
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1352;
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1353;
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1354;
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1355;
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1356;
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1357;
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1358;
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1359;
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1360;
  reg [31:0] _T_841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1361;
  reg [31:0] _T_841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1362;
  reg [31:0] _T_842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1363;
  reg [31:0] _T_842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1364;
  reg [31:0] _T_843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1365;
  reg [31:0] _T_843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1366;
  reg [31:0] _T_844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1367;
  reg [31:0] _T_844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1368;
  reg [31:0] _T_845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1369;
  reg [31:0] _T_845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1370;
  reg [31:0] _T_846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1371;
  reg [31:0] _T_846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1372;
  reg [31:0] _T_847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1373;
  reg [31:0] _T_847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1374;
  reg [31:0] _T_848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1375;
  reg [31:0] _T_848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1376;
  reg [31:0] _T_849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1377;
  reg [31:0] _T_849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1378;
  reg [31:0] _T_850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1379;
  reg [31:0] _T_850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1380;
  reg [31:0] _T_851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1381;
  reg [31:0] _T_851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1382;
  reg [31:0] _T_852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1383;
  reg [31:0] _T_852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1384;
  reg [31:0] _T_853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1385;
  reg [31:0] _T_853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1386;
  reg [31:0] _T_854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1387;
  reg [31:0] _T_854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1388;
  reg [31:0] _T_855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1389;
  reg [31:0] _T_855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1390;
  reg [31:0] _T_856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1391;
  reg [31:0] _T_856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1392;
  reg [31:0] _T_857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1393;
  reg [31:0] _T_857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1394;
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1395;
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1396;
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1397;
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1398;
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1399;
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1400;
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1401;
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1402;
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1403;
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1404;
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1405;
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1406;
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1407;
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1408;
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1409;
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1410;
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1411;
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1412;
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1413;
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1414;
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1415;
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1416;
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1417;
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1418;
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1419;
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1420;
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1421;
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1422;
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1423;
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1424;
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1425;
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1426;
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1427;
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1428;
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1429;
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1430;
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1431;
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1432;
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1433;
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1434;
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1435;
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1436;
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1437;
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1438;
  reg [31:0] _T_881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1439;
  reg [31:0] _T_881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1440;
  wire [31:0] _GEN_2402; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2403; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2404; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2405; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2406; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2407; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2408; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2409; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2410; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2411; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2412; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2413; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2414; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2415; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2418; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2419; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2420; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2421; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2422; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2423; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2424; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2425; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2426; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2427; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2428; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2429; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2430; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2431; // @[FFT.scala 35:12]
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1441;
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1442;
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1443;
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1444;
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1445;
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1446;
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1447;
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1448;
  reg [31:0] _T_890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1449;
  reg [31:0] _T_890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1450;
  reg [31:0] _T_891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1451;
  reg [31:0] _T_891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1452;
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1453;
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1454;
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1455;
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1456;
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1457;
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1458;
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1459;
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1460;
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1461;
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1462;
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1463;
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1464;
  reg [31:0] _T_898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1465;
  reg [31:0] _T_898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1466;
  reg [31:0] _T_899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1467;
  reg [31:0] _T_899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1468;
  reg [31:0] _T_900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1469;
  reg [31:0] _T_900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1470;
  reg [31:0] _T_901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1471;
  reg [31:0] _T_901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1472;
  reg [31:0] _T_903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1473;
  reg [31:0] _T_903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1474;
  reg [31:0] _T_904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1475;
  reg [31:0] _T_904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1476;
  reg [31:0] _T_905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1477;
  reg [31:0] _T_905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1478;
  reg [31:0] _T_906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1479;
  reg [31:0] _T_906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1480;
  reg [31:0] _T_907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1481;
  reg [31:0] _T_907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1482;
  reg [31:0] _T_908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1483;
  reg [31:0] _T_908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1484;
  reg [31:0] _T_909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1485;
  reg [31:0] _T_909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1486;
  reg [31:0] _T_910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1487;
  reg [31:0] _T_910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1488;
  wire [31:0] _GEN_2482; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2483; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2484; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2485; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2486; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2487; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2490; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2491; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2492; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2493; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2494; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2495; // @[FFT.scala 35:12]
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1489;
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1490;
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1491;
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1492;
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1493;
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1494;
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1495;
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1496;
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1497;
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1498;
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1499;
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1500;
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1501;
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1502;
  reg [31:0] _T_922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1503;
  reg [31:0] _T_922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1504;
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1505;
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1506;
  reg [31:0] _T_925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1507;
  reg [31:0] _T_925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1508;
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1509;
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1510;
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1511;
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1512;
  wire [31:0] _GEN_2522; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2523; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2526; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2527; // @[FFT.scala 35:12]
  reg [31:0] _T_932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1513;
  reg [31:0] _T_932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1514;
  reg [31:0] _T_933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1515;
  reg [31:0] _T_933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1516;
  reg [31:0] _T_934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1517;
  reg [31:0] _T_934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1518;
  reg [31:0] _T_935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1519;
  reg [31:0] _T_935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1520;
  reg [31:0] _T_937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1521;
  reg [31:0] _T_937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1522;
  reg [31:0] _T_938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1523;
  reg [31:0] _T_938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1524;
  reg [31:0] _T_943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1525;
  reg [31:0] _T_943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1526;
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1527;
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1528;
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1529;
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1530;
  reg [31:0] out1D1_re; // @[FFT.scala 58:23]
  reg [31:0] _RAND_1531;
  reg [31:0] out1D1_im; // @[FFT.scala 58:23]
  reg [31:0] _RAND_1532;
  reg [31:0] _T_947_re; // @[FFT.scala 62:22]
  reg [31:0] _RAND_1533;
  reg [31:0] _T_947_im; // @[FFT.scala 62:22]
  reg [31:0] _RAND_1534;
  reg [31:0] _T_948_re; // @[FFT.scala 63:22]
  reg [31:0] _RAND_1535;
  reg [31:0] _T_948_im; // @[FFT.scala 63:22]
  reg [31:0] _RAND_1536;
  reg  _T_949; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1537;
  reg  _T_950; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1538;
  reg  _T_951; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1539;
  reg  _T_952; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1540;
  reg  _T_953; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1541;
  reg  _T_954; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1542;
  reg  _T_955; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1543;
  reg  _T_956; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1544;
  reg  _T_957; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1545;
  reg  _T_958; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1546;
  reg  _T_959; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1547;
  reg  _T_960; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1548;
  reg  _T_961; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1549;
  reg  _T_962; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1550;
  reg  _T_963; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1551;
  reg  _T_964; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1552;
  reg  _T_965; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1553;
  reg  _T_966; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1554;
  reg  _T_967; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1555;
  reg  _T_968; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1556;
  reg  _T_969; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1557;
  reg  _T_970; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1558;
  reg  _T_971; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1559;
  reg  _T_972; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1560;
  reg  _T_973; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1561;
  reg  _T_974; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1562;
  reg  _T_975; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1563;
  reg  _T_976; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1564;
  reg  _T_977; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1565;
  reg  _T_978; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1566;
  reg  _T_979; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1567;
  reg  _T_980; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1568;
  reg  _T_981; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1569;
  reg  _T_982; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1570;
  reg  _T_983; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1571;
  reg  _T_984; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1572;
  reg  _T_985; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1573;
  reg  _T_986; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1574;
  reg  _T_987; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1575;
  reg  _T_988; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1576;
  reg  _T_989; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1577;
  reg  _T_990; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1578;
  reg  _T_991; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1579;
  reg  _T_992; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1580;
  reg  _T_993; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1581;
  reg  _T_994; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1582;
  reg  _T_995; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1583;
  reg  _T_996; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1584;
  reg  _T_997; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1585;
  reg  _T_998; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1586;
  reg  _T_999; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1587;
  reg  _T_1000; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1588;
  reg  _T_1001; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1589;
  reg  _T_1002; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1590;
  reg  _T_1003; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1591;
  reg  _T_1004; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1592;
  reg  _T_1005; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1593;
  reg  _T_1006; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1594;
  reg  _T_1007; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1595;
  reg  _T_1008; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1596;
  reg  _T_1009; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1597;
  reg  _T_1010; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1598;
  reg  _T_1011; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1599;
  reg  _T_1012; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1600;
  reg  _T_1013; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1601;
  reg  _T_1014; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1602;
  reg  _T_1015; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1603;
  reg  _T_1016; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1604;
  reg  _T_1017; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1605;
  reg  _T_1018; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1606;
  reg  _T_1019; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1607;
  reg  _T_1020; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1608;
  reg  _T_1021; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1609;
  reg  _T_1022; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1610;
  reg  _T_1023; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1611;
  reg  _T_1024; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1612;
  reg  _T_1025; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1613;
  reg  _T_1026; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1614;
  reg  _T_1027; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1615;
  reg  _T_1028; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1616;
  reg  _T_1029; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1617;
  reg  _T_1030; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1618;
  reg  _T_1031; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1619;
  reg  _T_1032; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1620;
  reg  _T_1033; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1621;
  reg  _T_1034; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1622;
  reg  _T_1035; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1623;
  reg  _T_1036; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1624;
  reg  _T_1037; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1625;
  reg  _T_1038; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1626;
  reg  _T_1039; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1627;
  reg  _T_1040; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1628;
  reg  _T_1041; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1629;
  reg  _T_1042; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1630;
  reg  _T_1043; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1631;
  reg  _T_1044; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1632;
  reg  _T_1045; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1633;
  reg  _T_1046; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1634;
  reg  _T_1047; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1635;
  reg  _T_1048; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1636;
  reg  _T_1049; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1637;
  reg  _T_1050; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1638;
  reg  _T_1051; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1639;
  reg  _T_1052; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1640;
  reg  _T_1053; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1641;
  reg  _T_1054; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1642;
  reg  _T_1055; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1643;
  reg  _T_1056; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1644;
  reg  _T_1057; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1645;
  reg  _T_1058; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1646;
  reg  _T_1059; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1647;
  reg  _T_1060; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1648;
  reg  _T_1061; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1649;
  reg  _T_1062; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1650;
  reg  _T_1063; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1651;
  reg  _T_1064; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1652;
  reg  _T_1065; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1653;
  reg  _T_1066; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1654;
  reg  _T_1067; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1655;
  reg  _T_1068; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1656;
  reg  _T_1069; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1657;
  reg  _T_1070; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1658;
  reg  _T_1071; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1659;
  reg  _T_1072; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1660;
  reg  _T_1073; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1661;
  reg  _T_1074; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1662;
  reg  _T_1075; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1663;
  reg  _T_1076; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1664;
  reg  _T_1077; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1665;
  reg  _T_1078; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1666;
  reg  _T_1079; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1667;
  reg  _T_1080; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1668;
  reg  _T_1081; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1669;
  reg  _T_1082; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1670;
  reg  _T_1083; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1671;
  reg  _T_1084; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1672;
  reg  _T_1085; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1673;
  reg  _T_1086; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1674;
  reg  _T_1087; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1675;
  reg  _T_1088; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1676;
  reg  _T_1089; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1677;
  reg  _T_1090; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1678;
  reg  _T_1091; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1679;
  reg  _T_1092; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1680;
  reg  _T_1093; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1681;
  reg  _T_1094; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1682;
  reg  _T_1095; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1683;
  reg  _T_1096; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1684;
  reg  _T_1097; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1685;
  reg  _T_1098; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1686;
  reg  _T_1099; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1687;
  reg  _T_1100; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1688;
  reg  _T_1101; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1689;
  reg  _T_1102; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1690;
  reg  _T_1103; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1691;
  reg  _T_1104; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1692;
  reg  _T_1105; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1693;
  reg  _T_1106; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1694;
  reg  _T_1107; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1695;
  reg  _T_1108; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1696;
  reg  _T_1109; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1697;
  reg  _T_1110; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1698;
  reg  _T_1111; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1699;
  reg  _T_1112; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1700;
  reg  _T_1113; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1701;
  reg  _T_1114; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1702;
  reg  _T_1115; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1703;
  reg  _T_1116; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1704;
  reg  _T_1117; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1705;
  reg  _T_1118; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1706;
  reg  _T_1119; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1707;
  reg  _T_1120; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1708;
  reg  _T_1121; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1709;
  reg  _T_1122; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1710;
  reg  _T_1123; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1711;
  reg  _T_1124; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1712;
  reg  _T_1125; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1713;
  reg  _T_1126; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1714;
  reg  _T_1127; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1715;
  reg  _T_1128; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1716;
  reg  _T_1129; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1717;
  reg  _T_1130; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1718;
  reg  _T_1131; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1719;
  reg  _T_1132; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1720;
  reg  _T_1133; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1721;
  reg  _T_1134; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1722;
  reg  _T_1135; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1723;
  reg  _T_1136; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1724;
  reg  _T_1137; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1725;
  reg  _T_1138; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1726;
  reg  _T_1139; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1727;
  reg  _T_1140; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1728;
  reg  _T_1141; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1729;
  reg  _T_1142; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1730;
  reg  _T_1143; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1731;
  reg  _T_1144; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1732;
  reg  _T_1145; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1733;
  reg  _T_1146; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1734;
  reg  _T_1147; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1735;
  reg  _T_1148; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1736;
  reg  _T_1149; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1737;
  reg  _T_1150; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1738;
  reg  _T_1151; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1739;
  reg  _T_1152; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1740;
  reg  _T_1153; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1741;
  reg  _T_1154; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1742;
  reg  _T_1155; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1743;
  reg  _T_1156; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1744;
  reg  _T_1157; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1745;
  reg  _T_1158; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1746;
  reg  _T_1159; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1747;
  reg  _T_1160; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1748;
  reg  _T_1161; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1749;
  reg  _T_1162; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1750;
  reg  _T_1163; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1751;
  reg  _T_1164; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1752;
  reg  _T_1165; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1753;
  reg  _T_1166; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1754;
  reg  _T_1167; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1755;
  reg  _T_1168; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1756;
  reg  _T_1169; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1757;
  reg  _T_1170; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1758;
  reg  _T_1171; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1759;
  reg  _T_1172; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1760;
  reg  _T_1173; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1761;
  reg  _T_1174; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1762;
  reg  _T_1175; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1763;
  reg  _T_1176; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1764;
  reg  _T_1177; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1765;
  reg  _T_1178; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1766;
  reg  _T_1179; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1767;
  reg  _T_1180; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1768;
  reg  _T_1181; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1769;
  reg  _T_1182; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1770;
  reg  _T_1183; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1771;
  reg  _T_1184; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1772;
  reg  _T_1185; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1773;
  reg  _T_1186; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1774;
  reg  _T_1187; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1775;
  reg  _T_1188; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1776;
  reg  _T_1189; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1777;
  reg  _T_1190; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1778;
  reg  _T_1191; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1779;
  reg  _T_1192; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1780;
  reg  _T_1193; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1781;
  reg  _T_1194; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1782;
  reg  _T_1195; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1783;
  reg  _T_1196; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1784;
  reg  _T_1197; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1785;
  reg  _T_1198; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1786;
  reg  _T_1199; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1787;
  reg  _T_1200; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1788;
  reg  _T_1201; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1789;
  reg  _T_1202; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1790;
  reg  _T_1203; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1791;
  reg  _T_1204; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1792;
  reg  _T_1205; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1793;
  reg  _T_1206; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1794;
  reg  _T_1207; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1795;
  reg  _T_1208; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1796;
  reg  _T_1209; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1797;
  reg  _T_1210; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1798;
  reg  _T_1211; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1799;
  reg  _T_1212; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1800;
  reg  _T_1213; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1801;
  reg  _T_1214; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1802;
  reg  _T_1215; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1803;
  reg  _T_1216; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1804;
  reg  _T_1217; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1805;
  reg  _T_1218; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1806;
  reg  _T_1219; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1807;
  reg  _T_1220; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1808;
  reg  _T_1221; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1809;
  reg  _T_1222; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1810;
  reg  _T_1223; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1811;
  reg  _T_1224; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1812;
  reg  _T_1225; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1813;
  reg  _T_1226; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1814;
  reg  _T_1227; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1815;
  reg  _T_1228; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1816;
  reg  _T_1229; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1817;
  reg  _T_1230; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1818;
  reg  _T_1231; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1819;
  reg  _T_1232; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1820;
  reg  _T_1233; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1821;
  reg  _T_1234; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1822;
  reg  _T_1235; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1823;
  reg  _T_1236; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1824;
  reg  _T_1237; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1825;
  reg  _T_1238; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1826;
  reg  _T_1239; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1827;
  reg  _T_1240; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1828;
  reg  _T_1241; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1829;
  reg  _T_1242; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1830;
  reg  _T_1243; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1831;
  reg  _T_1244; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1832;
  reg  _T_1245; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1833;
  reg  _T_1246; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1834;
  reg  _T_1247; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1835;
  reg  _T_1248; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1836;
  reg  _T_1249; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1837;
  reg  _T_1250; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1838;
  reg  _T_1251; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1839;
  reg  _T_1252; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1840;
  reg  _T_1253; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1841;
  reg  _T_1254; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1842;
  reg  _T_1255; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1843;
  reg  _T_1256; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1844;
  reg  _T_1257; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1845;
  reg  _T_1258; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1846;
  reg  _T_1259; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1847;
  reg  _T_1260; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1848;
  reg  _T_1261; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1849;
  reg  _T_1262; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1850;
  reg  _T_1263; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1851;
  reg  _T_1264; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1852;
  reg  _T_1265; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1853;
  reg  _T_1266; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1854;
  reg  _T_1267; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1855;
  reg  _T_1268; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1856;
  reg  _T_1269; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1857;
  reg  _T_1270; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1858;
  reg  _T_1271; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1859;
  reg  _T_1272; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1860;
  reg  _T_1273; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1861;
  reg  _T_1274; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1862;
  reg  _T_1275; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1863;
  reg  _T_1276; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1864;
  reg  _T_1277; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1865;
  reg  _T_1278; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1866;
  reg  _T_1279; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1867;
  reg  _T_1280; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1868;
  reg  _T_1281; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1869;
  reg  _T_1282; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1870;
  reg  _T_1283; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1871;
  reg  _T_1284; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1872;
  reg  _T_1285; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1873;
  reg  _T_1286; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1874;
  reg  _T_1287; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1875;
  reg  _T_1288; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1876;
  reg  _T_1289; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1877;
  reg  _T_1290; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1878;
  reg  _T_1291; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1879;
  reg  _T_1292; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1880;
  reg  _T_1293; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1881;
  reg  _T_1294; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1882;
  reg  _T_1295; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1883;
  reg  _T_1296; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1884;
  reg  _T_1297; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1885;
  reg  _T_1298; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1886;
  reg  _T_1299; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1887;
  reg  _T_1300; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1888;
  reg  _T_1301; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1889;
  reg  _T_1302; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1890;
  reg  _T_1303; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1891;
  reg  _T_1304; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1892;
  reg  _T_1305; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1893;
  reg  _T_1306; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1894;
  reg  _T_1307; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1895;
  reg  _T_1308; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1896;
  reg  _T_1309; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1897;
  reg  _T_1310; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1898;
  reg  _T_1311; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1899;
  reg  _T_1312; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1900;
  reg  _T_1313; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1901;
  reg  _T_1314; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1902;
  reg  _T_1315; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1903;
  reg  _T_1316; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1904;
  reg  _T_1317; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1905;
  reg  _T_1318; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1906;
  reg  _T_1319; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1907;
  reg  _T_1320; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1908;
  reg  _T_1321; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1909;
  reg  _T_1322; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1910;
  reg  _T_1323; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1911;
  reg  _T_1324; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1912;
  reg  _T_1325; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1913;
  reg  _T_1326; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1914;
  reg  _T_1327; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1915;
  reg  _T_1328; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1916;
  reg  _T_1329; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1917;
  reg  _T_1330; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1918;
  reg  _T_1331; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1919;
  reg  _T_1332; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1920;
  reg  _T_1333; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1921;
  reg  _T_1334; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1922;
  reg  _T_1335; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1923;
  reg  _T_1336; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1924;
  reg  _T_1337; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1925;
  reg  _T_1338; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1926;
  reg  _T_1339; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1927;
  reg  _T_1340; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1928;
  reg  _T_1341; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1929;
  reg  _T_1342; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1930;
  reg  _T_1343; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1931;
  reg  _T_1344; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1932;
  reg  _T_1345; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1933;
  reg  _T_1346; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1934;
  reg  _T_1347; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1935;
  reg  _T_1348; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1936;
  reg  _T_1349; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1937;
  reg  _T_1350; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1938;
  reg  _T_1351; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1939;
  reg  _T_1352; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1940;
  reg  _T_1353; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1941;
  reg  _T_1354; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1942;
  reg  _T_1355; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1943;
  reg  _T_1356; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1944;
  reg  _T_1357; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1945;
  reg  _T_1358; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1946;
  reg  _T_1359; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1947;
  reg  _T_1360; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1948;
  reg  _T_1361; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1949;
  reg  _T_1362; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1950;
  reg  _T_1363; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1951;
  reg  _T_1364; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1952;
  reg  _T_1365; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1953;
  reg  _T_1366; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1954;
  reg  _T_1367; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1955;
  reg  _T_1368; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1956;
  reg  _T_1369; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1957;
  reg  _T_1370; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1958;
  reg  _T_1371; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1959;
  reg  _T_1372; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1960;
  reg  _T_1373; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1961;
  reg  _T_1374; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1962;
  reg  _T_1375; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1963;
  reg  _T_1376; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1964;
  reg  _T_1377; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1965;
  reg  _T_1378; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1966;
  reg  _T_1379; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1967;
  reg  _T_1380; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1968;
  reg  _T_1381; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1969;
  reg  _T_1382; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1970;
  reg  _T_1383; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1971;
  reg  _T_1384; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1972;
  reg  _T_1385; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1973;
  reg  _T_1386; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1974;
  reg  _T_1387; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1975;
  reg  _T_1388; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1976;
  reg  _T_1389; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1977;
  reg  _T_1390; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1978;
  reg  _T_1391; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1979;
  reg  _T_1392; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1980;
  reg  _T_1393; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1981;
  reg  _T_1394; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1982;
  reg  _T_1395; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1983;
  reg  _T_1396; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1984;
  reg  _T_1397; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1985;
  reg  _T_1398; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1986;
  reg  _T_1399; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1987;
  reg  _T_1400; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1988;
  reg  _T_1401; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1989;
  reg  _T_1402; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1990;
  reg  _T_1403; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1991;
  reg  _T_1404; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1992;
  reg  _T_1405; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1993;
  reg  _T_1406; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1994;
  reg  _T_1407; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1995;
  reg  _T_1408; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1996;
  reg  _T_1409; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1997;
  reg  _T_1410; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1998;
  reg  _T_1411; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1999;
  reg  _T_1412; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2000;
  reg  _T_1413; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2001;
  reg  _T_1414; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2002;
  reg  _T_1415; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2003;
  reg  _T_1416; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2004;
  reg  _T_1417; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2005;
  reg  _T_1418; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2006;
  reg  _T_1419; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2007;
  reg  _T_1420; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2008;
  reg  _T_1421; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2009;
  reg  _T_1422; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2010;
  reg  _T_1423; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2011;
  reg  _T_1424; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2012;
  reg  _T_1425; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2013;
  reg  _T_1426; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2014;
  reg  _T_1427; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2015;
  reg  _T_1428; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2016;
  reg  _T_1429; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2017;
  reg  _T_1430; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2018;
  reg  _T_1431; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2019;
  reg  _T_1432; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2020;
  reg  _T_1433; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2021;
  reg  _T_1434; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2022;
  reg  _T_1435; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2023;
  reg  _T_1436; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2024;
  reg  _T_1437; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2025;
  reg  _T_1438; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2026;
  reg  _T_1439; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2027;
  reg  _T_1440; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2028;
  reg  _T_1441; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2029;
  reg  _T_1442; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2030;
  reg  _T_1443; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2031;
  reg  _T_1444; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2032;
  reg  _T_1445; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2033;
  reg  _T_1446; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2034;
  reg  _T_1447; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2035;
  reg  _T_1448; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2036;
  reg  _T_1449; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2037;
  reg  _T_1450; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2038;
  reg  _T_1451; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2039;
  reg  _T_1452; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2040;
  reg  _T_1453; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2041;
  reg  _T_1454; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2042;
  reg  _T_1455; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2043;
  reg  _T_1456; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2044;
  reg  _T_1457; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2045;
  reg  _T_1458; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2046;
  reg  _T_1459; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2047;
  reg  _T_1460; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2048;
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign _T_1 = cnt + 9'h1; // @[FFT.scala 42:16]
  assign _GEN_2 = 8'h1 == cnt[7:0] ? $signed(32'shfffb) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_3 = 8'h2 == cnt[7:0] ? $signed(32'shffec) : $signed(_GEN_2); // @[FFT.scala 34:12]
  assign _GEN_4 = 8'h3 == cnt[7:0] ? $signed(32'shffd4) : $signed(_GEN_3); // @[FFT.scala 34:12]
  assign _GEN_5 = 8'h4 == cnt[7:0] ? $signed(32'shffb1) : $signed(_GEN_4); // @[FFT.scala 34:12]
  assign _GEN_6 = 8'h5 == cnt[7:0] ? $signed(32'shff85) : $signed(_GEN_5); // @[FFT.scala 34:12]
  assign _GEN_7 = 8'h6 == cnt[7:0] ? $signed(32'shff4e) : $signed(_GEN_6); // @[FFT.scala 34:12]
  assign _GEN_8 = 8'h7 == cnt[7:0] ? $signed(32'shff0e) : $signed(_GEN_7); // @[FFT.scala 34:12]
  assign _GEN_9 = 8'h8 == cnt[7:0] ? $signed(32'shfec4) : $signed(_GEN_8); // @[FFT.scala 34:12]
  assign _GEN_10 = 8'h9 == cnt[7:0] ? $signed(32'shfe71) : $signed(_GEN_9); // @[FFT.scala 34:12]
  assign _GEN_11 = 8'ha == cnt[7:0] ? $signed(32'shfe13) : $signed(_GEN_10); // @[FFT.scala 34:12]
  assign _GEN_12 = 8'hb == cnt[7:0] ? $signed(32'shfdac) : $signed(_GEN_11); // @[FFT.scala 34:12]
  assign _GEN_13 = 8'hc == cnt[7:0] ? $signed(32'shfd3b) : $signed(_GEN_12); // @[FFT.scala 34:12]
  assign _GEN_14 = 8'hd == cnt[7:0] ? $signed(32'shfcc0) : $signed(_GEN_13); // @[FFT.scala 34:12]
  assign _GEN_15 = 8'he == cnt[7:0] ? $signed(32'shfc3b) : $signed(_GEN_14); // @[FFT.scala 34:12]
  assign _GEN_16 = 8'hf == cnt[7:0] ? $signed(32'shfbad) : $signed(_GEN_15); // @[FFT.scala 34:12]
  assign _GEN_17 = 8'h10 == cnt[7:0] ? $signed(32'shfb15) : $signed(_GEN_16); // @[FFT.scala 34:12]
  assign _GEN_18 = 8'h11 == cnt[7:0] ? $signed(32'shfa73) : $signed(_GEN_17); // @[FFT.scala 34:12]
  assign _GEN_19 = 8'h12 == cnt[7:0] ? $signed(32'shf9c8) : $signed(_GEN_18); // @[FFT.scala 34:12]
  assign _GEN_20 = 8'h13 == cnt[7:0] ? $signed(32'shf913) : $signed(_GEN_19); // @[FFT.scala 34:12]
  assign _GEN_21 = 8'h14 == cnt[7:0] ? $signed(32'shf854) : $signed(_GEN_20); // @[FFT.scala 34:12]
  assign _GEN_22 = 8'h15 == cnt[7:0] ? $signed(32'shf78c) : $signed(_GEN_21); // @[FFT.scala 34:12]
  assign _GEN_23 = 8'h16 == cnt[7:0] ? $signed(32'shf6ba) : $signed(_GEN_22); // @[FFT.scala 34:12]
  assign _GEN_24 = 8'h17 == cnt[7:0] ? $signed(32'shf5df) : $signed(_GEN_23); // @[FFT.scala 34:12]
  assign _GEN_25 = 8'h18 == cnt[7:0] ? $signed(32'shf4fa) : $signed(_GEN_24); // @[FFT.scala 34:12]
  assign _GEN_26 = 8'h19 == cnt[7:0] ? $signed(32'shf40c) : $signed(_GEN_25); // @[FFT.scala 34:12]
  assign _GEN_27 = 8'h1a == cnt[7:0] ? $signed(32'shf314) : $signed(_GEN_26); // @[FFT.scala 34:12]
  assign _GEN_28 = 8'h1b == cnt[7:0] ? $signed(32'shf213) : $signed(_GEN_27); // @[FFT.scala 34:12]
  assign _GEN_29 = 8'h1c == cnt[7:0] ? $signed(32'shf109) : $signed(_GEN_28); // @[FFT.scala 34:12]
  assign _GEN_30 = 8'h1d == cnt[7:0] ? $signed(32'sheff5) : $signed(_GEN_29); // @[FFT.scala 34:12]
  assign _GEN_31 = 8'h1e == cnt[7:0] ? $signed(32'sheed9) : $signed(_GEN_30); // @[FFT.scala 34:12]
  assign _GEN_32 = 8'h1f == cnt[7:0] ? $signed(32'shedb3) : $signed(_GEN_31); // @[FFT.scala 34:12]
  assign _GEN_33 = 8'h20 == cnt[7:0] ? $signed(32'shec83) : $signed(_GEN_32); // @[FFT.scala 34:12]
  assign _GEN_34 = 8'h21 == cnt[7:0] ? $signed(32'sheb4b) : $signed(_GEN_33); // @[FFT.scala 34:12]
  assign _GEN_35 = 8'h22 == cnt[7:0] ? $signed(32'shea0a) : $signed(_GEN_34); // @[FFT.scala 34:12]
  assign _GEN_36 = 8'h23 == cnt[7:0] ? $signed(32'she8bf) : $signed(_GEN_35); // @[FFT.scala 34:12]
  assign _GEN_37 = 8'h24 == cnt[7:0] ? $signed(32'she76c) : $signed(_GEN_36); // @[FFT.scala 34:12]
  assign _GEN_38 = 8'h25 == cnt[7:0] ? $signed(32'she610) : $signed(_GEN_37); // @[FFT.scala 34:12]
  assign _GEN_39 = 8'h26 == cnt[7:0] ? $signed(32'she4aa) : $signed(_GEN_38); // @[FFT.scala 34:12]
  assign _GEN_40 = 8'h27 == cnt[7:0] ? $signed(32'she33c) : $signed(_GEN_39); // @[FFT.scala 34:12]
  assign _GEN_41 = 8'h28 == cnt[7:0] ? $signed(32'she1c6) : $signed(_GEN_40); // @[FFT.scala 34:12]
  assign _GEN_42 = 8'h29 == cnt[7:0] ? $signed(32'she046) : $signed(_GEN_41); // @[FFT.scala 34:12]
  assign _GEN_43 = 8'h2a == cnt[7:0] ? $signed(32'shdebe) : $signed(_GEN_42); // @[FFT.scala 34:12]
  assign _GEN_44 = 8'h2b == cnt[7:0] ? $signed(32'shdd2d) : $signed(_GEN_43); // @[FFT.scala 34:12]
  assign _GEN_45 = 8'h2c == cnt[7:0] ? $signed(32'shdb94) : $signed(_GEN_44); // @[FFT.scala 34:12]
  assign _GEN_46 = 8'h2d == cnt[7:0] ? $signed(32'shd9f2) : $signed(_GEN_45); // @[FFT.scala 34:12]
  assign _GEN_47 = 8'h2e == cnt[7:0] ? $signed(32'shd848) : $signed(_GEN_46); // @[FFT.scala 34:12]
  assign _GEN_48 = 8'h2f == cnt[7:0] ? $signed(32'shd696) : $signed(_GEN_47); // @[FFT.scala 34:12]
  assign _GEN_49 = 8'h30 == cnt[7:0] ? $signed(32'shd4db) : $signed(_GEN_48); // @[FFT.scala 34:12]
  assign _GEN_50 = 8'h31 == cnt[7:0] ? $signed(32'shd318) : $signed(_GEN_49); // @[FFT.scala 34:12]
  assign _GEN_51 = 8'h32 == cnt[7:0] ? $signed(32'shd14d) : $signed(_GEN_50); // @[FFT.scala 34:12]
  assign _GEN_52 = 8'h33 == cnt[7:0] ? $signed(32'shcf7a) : $signed(_GEN_51); // @[FFT.scala 34:12]
  assign _GEN_53 = 8'h34 == cnt[7:0] ? $signed(32'shcd9f) : $signed(_GEN_52); // @[FFT.scala 34:12]
  assign _GEN_54 = 8'h35 == cnt[7:0] ? $signed(32'shcbbc) : $signed(_GEN_53); // @[FFT.scala 34:12]
  assign _GEN_55 = 8'h36 == cnt[7:0] ? $signed(32'shc9d1) : $signed(_GEN_54); // @[FFT.scala 34:12]
  assign _GEN_56 = 8'h37 == cnt[7:0] ? $signed(32'shc7de) : $signed(_GEN_55); // @[FFT.scala 34:12]
  assign _GEN_57 = 8'h38 == cnt[7:0] ? $signed(32'shc5e4) : $signed(_GEN_56); // @[FFT.scala 34:12]
  assign _GEN_58 = 8'h39 == cnt[7:0] ? $signed(32'shc3e2) : $signed(_GEN_57); // @[FFT.scala 34:12]
  assign _GEN_59 = 8'h3a == cnt[7:0] ? $signed(32'shc1d8) : $signed(_GEN_58); // @[FFT.scala 34:12]
  assign _GEN_60 = 8'h3b == cnt[7:0] ? $signed(32'shbfc7) : $signed(_GEN_59); // @[FFT.scala 34:12]
  assign _GEN_61 = 8'h3c == cnt[7:0] ? $signed(32'shbdaf) : $signed(_GEN_60); // @[FFT.scala 34:12]
  assign _GEN_62 = 8'h3d == cnt[7:0] ? $signed(32'shbb8f) : $signed(_GEN_61); // @[FFT.scala 34:12]
  assign _GEN_63 = 8'h3e == cnt[7:0] ? $signed(32'shb968) : $signed(_GEN_62); // @[FFT.scala 34:12]
  assign _GEN_64 = 8'h3f == cnt[7:0] ? $signed(32'shb73a) : $signed(_GEN_63); // @[FFT.scala 34:12]
  assign _GEN_65 = 8'h40 == cnt[7:0] ? $signed(32'shb505) : $signed(_GEN_64); // @[FFT.scala 34:12]
  assign _GEN_66 = 8'h41 == cnt[7:0] ? $signed(32'shb2c9) : $signed(_GEN_65); // @[FFT.scala 34:12]
  assign _GEN_67 = 8'h42 == cnt[7:0] ? $signed(32'shb086) : $signed(_GEN_66); // @[FFT.scala 34:12]
  assign _GEN_68 = 8'h43 == cnt[7:0] ? $signed(32'shae3c) : $signed(_GEN_67); // @[FFT.scala 34:12]
  assign _GEN_69 = 8'h44 == cnt[7:0] ? $signed(32'shabeb) : $signed(_GEN_68); // @[FFT.scala 34:12]
  assign _GEN_70 = 8'h45 == cnt[7:0] ? $signed(32'sha994) : $signed(_GEN_69); // @[FFT.scala 34:12]
  assign _GEN_71 = 8'h46 == cnt[7:0] ? $signed(32'sha736) : $signed(_GEN_70); // @[FFT.scala 34:12]
  assign _GEN_72 = 8'h47 == cnt[7:0] ? $signed(32'sha4d2) : $signed(_GEN_71); // @[FFT.scala 34:12]
  assign _GEN_73 = 8'h48 == cnt[7:0] ? $signed(32'sha268) : $signed(_GEN_72); // @[FFT.scala 34:12]
  assign _GEN_74 = 8'h49 == cnt[7:0] ? $signed(32'sh9ff7) : $signed(_GEN_73); // @[FFT.scala 34:12]
  assign _GEN_75 = 8'h4a == cnt[7:0] ? $signed(32'sh9d80) : $signed(_GEN_74); // @[FFT.scala 34:12]
  assign _GEN_76 = 8'h4b == cnt[7:0] ? $signed(32'sh9b03) : $signed(_GEN_75); // @[FFT.scala 34:12]
  assign _GEN_77 = 8'h4c == cnt[7:0] ? $signed(32'sh9880) : $signed(_GEN_76); // @[FFT.scala 34:12]
  assign _GEN_78 = 8'h4d == cnt[7:0] ? $signed(32'sh95f7) : $signed(_GEN_77); // @[FFT.scala 34:12]
  assign _GEN_79 = 8'h4e == cnt[7:0] ? $signed(32'sh9368) : $signed(_GEN_78); // @[FFT.scala 34:12]
  assign _GEN_80 = 8'h4f == cnt[7:0] ? $signed(32'sh90d4) : $signed(_GEN_79); // @[FFT.scala 34:12]
  assign _GEN_81 = 8'h50 == cnt[7:0] ? $signed(32'sh8e3a) : $signed(_GEN_80); // @[FFT.scala 34:12]
  assign _GEN_82 = 8'h51 == cnt[7:0] ? $signed(32'sh8b9a) : $signed(_GEN_81); // @[FFT.scala 34:12]
  assign _GEN_83 = 8'h52 == cnt[7:0] ? $signed(32'sh88f6) : $signed(_GEN_82); // @[FFT.scala 34:12]
  assign _GEN_84 = 8'h53 == cnt[7:0] ? $signed(32'sh864c) : $signed(_GEN_83); // @[FFT.scala 34:12]
  assign _GEN_85 = 8'h54 == cnt[7:0] ? $signed(32'sh839c) : $signed(_GEN_84); // @[FFT.scala 34:12]
  assign _GEN_86 = 8'h55 == cnt[7:0] ? $signed(32'sh80e8) : $signed(_GEN_85); // @[FFT.scala 34:12]
  assign _GEN_87 = 8'h56 == cnt[7:0] ? $signed(32'sh7e2f) : $signed(_GEN_86); // @[FFT.scala 34:12]
  assign _GEN_88 = 8'h57 == cnt[7:0] ? $signed(32'sh7b70) : $signed(_GEN_87); // @[FFT.scala 34:12]
  assign _GEN_89 = 8'h58 == cnt[7:0] ? $signed(32'sh78ad) : $signed(_GEN_88); // @[FFT.scala 34:12]
  assign _GEN_90 = 8'h59 == cnt[7:0] ? $signed(32'sh75e6) : $signed(_GEN_89); // @[FFT.scala 34:12]
  assign _GEN_91 = 8'h5a == cnt[7:0] ? $signed(32'sh731a) : $signed(_GEN_90); // @[FFT.scala 34:12]
  assign _GEN_92 = 8'h5b == cnt[7:0] ? $signed(32'sh7049) : $signed(_GEN_91); // @[FFT.scala 34:12]
  assign _GEN_93 = 8'h5c == cnt[7:0] ? $signed(32'sh6d74) : $signed(_GEN_92); // @[FFT.scala 34:12]
  assign _GEN_94 = 8'h5d == cnt[7:0] ? $signed(32'sh6a9b) : $signed(_GEN_93); // @[FFT.scala 34:12]
  assign _GEN_95 = 8'h5e == cnt[7:0] ? $signed(32'sh67be) : $signed(_GEN_94); // @[FFT.scala 34:12]
  assign _GEN_96 = 8'h5f == cnt[7:0] ? $signed(32'sh64dd) : $signed(_GEN_95); // @[FFT.scala 34:12]
  assign _GEN_97 = 8'h60 == cnt[7:0] ? $signed(32'sh61f8) : $signed(_GEN_96); // @[FFT.scala 34:12]
  assign _GEN_98 = 8'h61 == cnt[7:0] ? $signed(32'sh5f0f) : $signed(_GEN_97); // @[FFT.scala 34:12]
  assign _GEN_99 = 8'h62 == cnt[7:0] ? $signed(32'sh5c22) : $signed(_GEN_98); // @[FFT.scala 34:12]
  assign _GEN_100 = 8'h63 == cnt[7:0] ? $signed(32'sh5932) : $signed(_GEN_99); // @[FFT.scala 34:12]
  assign _GEN_101 = 8'h64 == cnt[7:0] ? $signed(32'sh563e) : $signed(_GEN_100); // @[FFT.scala 34:12]
  assign _GEN_102 = 8'h65 == cnt[7:0] ? $signed(32'sh5348) : $signed(_GEN_101); // @[FFT.scala 34:12]
  assign _GEN_103 = 8'h66 == cnt[7:0] ? $signed(32'sh504d) : $signed(_GEN_102); // @[FFT.scala 34:12]
  assign _GEN_104 = 8'h67 == cnt[7:0] ? $signed(32'sh4d50) : $signed(_GEN_103); // @[FFT.scala 34:12]
  assign _GEN_105 = 8'h68 == cnt[7:0] ? $signed(32'sh4a50) : $signed(_GEN_104); // @[FFT.scala 34:12]
  assign _GEN_106 = 8'h69 == cnt[7:0] ? $signed(32'sh474d) : $signed(_GEN_105); // @[FFT.scala 34:12]
  assign _GEN_107 = 8'h6a == cnt[7:0] ? $signed(32'sh4447) : $signed(_GEN_106); // @[FFT.scala 34:12]
  assign _GEN_108 = 8'h6b == cnt[7:0] ? $signed(32'sh413f) : $signed(_GEN_107); // @[FFT.scala 34:12]
  assign _GEN_109 = 8'h6c == cnt[7:0] ? $signed(32'sh3e34) : $signed(_GEN_108); // @[FFT.scala 34:12]
  assign _GEN_110 = 8'h6d == cnt[7:0] ? $signed(32'sh3b27) : $signed(_GEN_109); // @[FFT.scala 34:12]
  assign _GEN_111 = 8'h6e == cnt[7:0] ? $signed(32'sh3817) : $signed(_GEN_110); // @[FFT.scala 34:12]
  assign _GEN_112 = 8'h6f == cnt[7:0] ? $signed(32'sh3505) : $signed(_GEN_111); // @[FFT.scala 34:12]
  assign _GEN_113 = 8'h70 == cnt[7:0] ? $signed(32'sh31f1) : $signed(_GEN_112); // @[FFT.scala 34:12]
  assign _GEN_114 = 8'h71 == cnt[7:0] ? $signed(32'sh2edc) : $signed(_GEN_113); // @[FFT.scala 34:12]
  assign _GEN_115 = 8'h72 == cnt[7:0] ? $signed(32'sh2bc4) : $signed(_GEN_114); // @[FFT.scala 34:12]
  assign _GEN_116 = 8'h73 == cnt[7:0] ? $signed(32'sh28ab) : $signed(_GEN_115); // @[FFT.scala 34:12]
  assign _GEN_117 = 8'h74 == cnt[7:0] ? $signed(32'sh2590) : $signed(_GEN_116); // @[FFT.scala 34:12]
  assign _GEN_118 = 8'h75 == cnt[7:0] ? $signed(32'sh2274) : $signed(_GEN_117); // @[FFT.scala 34:12]
  assign _GEN_119 = 8'h76 == cnt[7:0] ? $signed(32'sh1f56) : $signed(_GEN_118); // @[FFT.scala 34:12]
  assign _GEN_120 = 8'h77 == cnt[7:0] ? $signed(32'sh1c38) : $signed(_GEN_119); // @[FFT.scala 34:12]
  assign _GEN_121 = 8'h78 == cnt[7:0] ? $signed(32'sh1918) : $signed(_GEN_120); // @[FFT.scala 34:12]
  assign _GEN_122 = 8'h79 == cnt[7:0] ? $signed(32'sh15f7) : $signed(_GEN_121); // @[FFT.scala 34:12]
  assign _GEN_123 = 8'h7a == cnt[7:0] ? $signed(32'sh12d5) : $signed(_GEN_122); // @[FFT.scala 34:12]
  assign _GEN_124 = 8'h7b == cnt[7:0] ? $signed(32'shfb3) : $signed(_GEN_123); // @[FFT.scala 34:12]
  assign _GEN_125 = 8'h7c == cnt[7:0] ? $signed(32'shc90) : $signed(_GEN_124); // @[FFT.scala 34:12]
  assign _GEN_126 = 8'h7d == cnt[7:0] ? $signed(32'sh96c) : $signed(_GEN_125); // @[FFT.scala 34:12]
  assign _GEN_127 = 8'h7e == cnt[7:0] ? $signed(32'sh648) : $signed(_GEN_126); // @[FFT.scala 34:12]
  assign _GEN_128 = 8'h7f == cnt[7:0] ? $signed(32'sh324) : $signed(_GEN_127); // @[FFT.scala 34:12]
  assign _GEN_129 = 8'h80 == cnt[7:0] ? $signed(32'sh0) : $signed(_GEN_128); // @[FFT.scala 34:12]
  assign _GEN_130 = 8'h81 == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_129); // @[FFT.scala 34:12]
  assign _GEN_131 = 8'h82 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_130); // @[FFT.scala 34:12]
  assign _GEN_132 = 8'h83 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_131); // @[FFT.scala 34:12]
  assign _GEN_133 = 8'h84 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_132); // @[FFT.scala 34:12]
  assign _GEN_134 = 8'h85 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_133); // @[FFT.scala 34:12]
  assign _GEN_135 = 8'h86 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_134); // @[FFT.scala 34:12]
  assign _GEN_136 = 8'h87 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_135); // @[FFT.scala 34:12]
  assign _GEN_137 = 8'h88 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_136); // @[FFT.scala 34:12]
  assign _GEN_138 = 8'h89 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_137); // @[FFT.scala 34:12]
  assign _GEN_139 = 8'h8a == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_138); // @[FFT.scala 34:12]
  assign _GEN_140 = 8'h8b == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_139); // @[FFT.scala 34:12]
  assign _GEN_141 = 8'h8c == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_140); // @[FFT.scala 34:12]
  assign _GEN_142 = 8'h8d == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_141); // @[FFT.scala 34:12]
  assign _GEN_143 = 8'h8e == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_142); // @[FFT.scala 34:12]
  assign _GEN_144 = 8'h8f == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_143); // @[FFT.scala 34:12]
  assign _GEN_145 = 8'h90 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_144); // @[FFT.scala 34:12]
  assign _GEN_146 = 8'h91 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_145); // @[FFT.scala 34:12]
  assign _GEN_147 = 8'h92 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_146); // @[FFT.scala 34:12]
  assign _GEN_148 = 8'h93 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_147); // @[FFT.scala 34:12]
  assign _GEN_149 = 8'h94 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_148); // @[FFT.scala 34:12]
  assign _GEN_150 = 8'h95 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_149); // @[FFT.scala 34:12]
  assign _GEN_151 = 8'h96 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_150); // @[FFT.scala 34:12]
  assign _GEN_152 = 8'h97 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_151); // @[FFT.scala 34:12]
  assign _GEN_153 = 8'h98 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_152); // @[FFT.scala 34:12]
  assign _GEN_154 = 8'h99 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_153); // @[FFT.scala 34:12]
  assign _GEN_155 = 8'h9a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_154); // @[FFT.scala 34:12]
  assign _GEN_156 = 8'h9b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_155); // @[FFT.scala 34:12]
  assign _GEN_157 = 8'h9c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_156); // @[FFT.scala 34:12]
  assign _GEN_158 = 8'h9d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_157); // @[FFT.scala 34:12]
  assign _GEN_159 = 8'h9e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_158); // @[FFT.scala 34:12]
  assign _GEN_160 = 8'h9f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_159); // @[FFT.scala 34:12]
  assign _GEN_161 = 8'ha0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_160); // @[FFT.scala 34:12]
  assign _GEN_162 = 8'ha1 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_161); // @[FFT.scala 34:12]
  assign _GEN_163 = 8'ha2 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_162); // @[FFT.scala 34:12]
  assign _GEN_164 = 8'ha3 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_163); // @[FFT.scala 34:12]
  assign _GEN_165 = 8'ha4 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_164); // @[FFT.scala 34:12]
  assign _GEN_166 = 8'ha5 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_165); // @[FFT.scala 34:12]
  assign _GEN_167 = 8'ha6 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_166); // @[FFT.scala 34:12]
  assign _GEN_168 = 8'ha7 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_167); // @[FFT.scala 34:12]
  assign _GEN_169 = 8'ha8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_168); // @[FFT.scala 34:12]
  assign _GEN_170 = 8'ha9 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_169); // @[FFT.scala 34:12]
  assign _GEN_171 = 8'haa == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_170); // @[FFT.scala 34:12]
  assign _GEN_172 = 8'hab == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_171); // @[FFT.scala 34:12]
  assign _GEN_173 = 8'hac == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_172); // @[FFT.scala 34:12]
  assign _GEN_174 = 8'had == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_173); // @[FFT.scala 34:12]
  assign _GEN_175 = 8'hae == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_174); // @[FFT.scala 34:12]
  assign _GEN_176 = 8'haf == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_175); // @[FFT.scala 34:12]
  assign _GEN_177 = 8'hb0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_176); // @[FFT.scala 34:12]
  assign _GEN_178 = 8'hb1 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_177); // @[FFT.scala 34:12]
  assign _GEN_179 = 8'hb2 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_178); // @[FFT.scala 34:12]
  assign _GEN_180 = 8'hb3 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_179); // @[FFT.scala 34:12]
  assign _GEN_181 = 8'hb4 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_180); // @[FFT.scala 34:12]
  assign _GEN_182 = 8'hb5 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_181); // @[FFT.scala 34:12]
  assign _GEN_183 = 8'hb6 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_182); // @[FFT.scala 34:12]
  assign _GEN_184 = 8'hb7 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_183); // @[FFT.scala 34:12]
  assign _GEN_185 = 8'hb8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_184); // @[FFT.scala 34:12]
  assign _GEN_186 = 8'hb9 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_185); // @[FFT.scala 34:12]
  assign _GEN_187 = 8'hba == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_186); // @[FFT.scala 34:12]
  assign _GEN_188 = 8'hbb == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_187); // @[FFT.scala 34:12]
  assign _GEN_189 = 8'hbc == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_188); // @[FFT.scala 34:12]
  assign _GEN_190 = 8'hbd == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_189); // @[FFT.scala 34:12]
  assign _GEN_191 = 8'hbe == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_190); // @[FFT.scala 34:12]
  assign _GEN_192 = 8'hbf == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_191); // @[FFT.scala 34:12]
  assign _GEN_193 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_192); // @[FFT.scala 34:12]
  assign _GEN_194 = 8'hc1 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_193); // @[FFT.scala 34:12]
  assign _GEN_195 = 8'hc2 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_194); // @[FFT.scala 34:12]
  assign _GEN_196 = 8'hc3 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_195); // @[FFT.scala 34:12]
  assign _GEN_197 = 8'hc4 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_196); // @[FFT.scala 34:12]
  assign _GEN_198 = 8'hc5 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_197); // @[FFT.scala 34:12]
  assign _GEN_199 = 8'hc6 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_198); // @[FFT.scala 34:12]
  assign _GEN_200 = 8'hc7 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_199); // @[FFT.scala 34:12]
  assign _GEN_201 = 8'hc8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_200); // @[FFT.scala 34:12]
  assign _GEN_202 = 8'hc9 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_201); // @[FFT.scala 34:12]
  assign _GEN_203 = 8'hca == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_202); // @[FFT.scala 34:12]
  assign _GEN_204 = 8'hcb == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_203); // @[FFT.scala 34:12]
  assign _GEN_205 = 8'hcc == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_204); // @[FFT.scala 34:12]
  assign _GEN_206 = 8'hcd == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_205); // @[FFT.scala 34:12]
  assign _GEN_207 = 8'hce == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_206); // @[FFT.scala 34:12]
  assign _GEN_208 = 8'hcf == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_207); // @[FFT.scala 34:12]
  assign _GEN_209 = 8'hd0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_208); // @[FFT.scala 34:12]
  assign _GEN_210 = 8'hd1 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_209); // @[FFT.scala 34:12]
  assign _GEN_211 = 8'hd2 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_210); // @[FFT.scala 34:12]
  assign _GEN_212 = 8'hd3 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_211); // @[FFT.scala 34:12]
  assign _GEN_213 = 8'hd4 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_212); // @[FFT.scala 34:12]
  assign _GEN_214 = 8'hd5 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_213); // @[FFT.scala 34:12]
  assign _GEN_215 = 8'hd6 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_214); // @[FFT.scala 34:12]
  assign _GEN_216 = 8'hd7 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_215); // @[FFT.scala 34:12]
  assign _GEN_217 = 8'hd8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_216); // @[FFT.scala 34:12]
  assign _GEN_218 = 8'hd9 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_217); // @[FFT.scala 34:12]
  assign _GEN_219 = 8'hda == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_218); // @[FFT.scala 34:12]
  assign _GEN_220 = 8'hdb == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_219); // @[FFT.scala 34:12]
  assign _GEN_221 = 8'hdc == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_220); // @[FFT.scala 34:12]
  assign _GEN_222 = 8'hdd == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_221); // @[FFT.scala 34:12]
  assign _GEN_223 = 8'hde == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_222); // @[FFT.scala 34:12]
  assign _GEN_224 = 8'hdf == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_223); // @[FFT.scala 34:12]
  assign _GEN_225 = 8'he0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_224); // @[FFT.scala 34:12]
  assign _GEN_226 = 8'he1 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_225); // @[FFT.scala 34:12]
  assign _GEN_227 = 8'he2 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_226); // @[FFT.scala 34:12]
  assign _GEN_228 = 8'he3 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_227); // @[FFT.scala 34:12]
  assign _GEN_229 = 8'he4 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_228); // @[FFT.scala 34:12]
  assign _GEN_230 = 8'he5 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_229); // @[FFT.scala 34:12]
  assign _GEN_231 = 8'he6 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_230); // @[FFT.scala 34:12]
  assign _GEN_232 = 8'he7 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_231); // @[FFT.scala 34:12]
  assign _GEN_233 = 8'he8 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_232); // @[FFT.scala 34:12]
  assign _GEN_234 = 8'he9 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_233); // @[FFT.scala 34:12]
  assign _GEN_235 = 8'hea == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_234); // @[FFT.scala 34:12]
  assign _GEN_236 = 8'heb == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_235); // @[FFT.scala 34:12]
  assign _GEN_237 = 8'hec == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_236); // @[FFT.scala 34:12]
  assign _GEN_238 = 8'hed == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_237); // @[FFT.scala 34:12]
  assign _GEN_239 = 8'hee == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_238); // @[FFT.scala 34:12]
  assign _GEN_240 = 8'hef == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_239); // @[FFT.scala 34:12]
  assign _GEN_241 = 8'hf0 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_240); // @[FFT.scala 34:12]
  assign _GEN_242 = 8'hf1 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_241); // @[FFT.scala 34:12]
  assign _GEN_243 = 8'hf2 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_242); // @[FFT.scala 34:12]
  assign _GEN_244 = 8'hf3 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_243); // @[FFT.scala 34:12]
  assign _GEN_245 = 8'hf4 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_244); // @[FFT.scala 34:12]
  assign _GEN_246 = 8'hf5 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_245); // @[FFT.scala 34:12]
  assign _GEN_247 = 8'hf6 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_246); // @[FFT.scala 34:12]
  assign _GEN_248 = 8'hf7 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_247); // @[FFT.scala 34:12]
  assign _GEN_249 = 8'hf8 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_248); // @[FFT.scala 34:12]
  assign _GEN_250 = 8'hf9 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_249); // @[FFT.scala 34:12]
  assign _GEN_251 = 8'hfa == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_250); // @[FFT.scala 34:12]
  assign _GEN_252 = 8'hfb == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_251); // @[FFT.scala 34:12]
  assign _GEN_253 = 8'hfc == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_252); // @[FFT.scala 34:12]
  assign _GEN_254 = 8'hfd == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_253); // @[FFT.scala 34:12]
  assign _GEN_255 = 8'hfe == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_254); // @[FFT.scala 34:12]
  assign _GEN_258 = 8'h1 == cnt[7:0] ? $signed(-32'sh324) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_259 = 8'h2 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_258); // @[FFT.scala 35:12]
  assign _GEN_260 = 8'h3 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_259); // @[FFT.scala 35:12]
  assign _GEN_261 = 8'h4 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_260); // @[FFT.scala 35:12]
  assign _GEN_262 = 8'h5 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_261); // @[FFT.scala 35:12]
  assign _GEN_263 = 8'h6 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_262); // @[FFT.scala 35:12]
  assign _GEN_264 = 8'h7 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_263); // @[FFT.scala 35:12]
  assign _GEN_265 = 8'h8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_264); // @[FFT.scala 35:12]
  assign _GEN_266 = 8'h9 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_265); // @[FFT.scala 35:12]
  assign _GEN_267 = 8'ha == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_266); // @[FFT.scala 35:12]
  assign _GEN_268 = 8'hb == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_267); // @[FFT.scala 35:12]
  assign _GEN_269 = 8'hc == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_268); // @[FFT.scala 35:12]
  assign _GEN_270 = 8'hd == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_269); // @[FFT.scala 35:12]
  assign _GEN_271 = 8'he == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_270); // @[FFT.scala 35:12]
  assign _GEN_272 = 8'hf == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_271); // @[FFT.scala 35:12]
  assign _GEN_273 = 8'h10 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_272); // @[FFT.scala 35:12]
  assign _GEN_274 = 8'h11 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_273); // @[FFT.scala 35:12]
  assign _GEN_275 = 8'h12 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_274); // @[FFT.scala 35:12]
  assign _GEN_276 = 8'h13 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_275); // @[FFT.scala 35:12]
  assign _GEN_277 = 8'h14 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_276); // @[FFT.scala 35:12]
  assign _GEN_278 = 8'h15 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_277); // @[FFT.scala 35:12]
  assign _GEN_279 = 8'h16 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_278); // @[FFT.scala 35:12]
  assign _GEN_280 = 8'h17 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_279); // @[FFT.scala 35:12]
  assign _GEN_281 = 8'h18 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_280); // @[FFT.scala 35:12]
  assign _GEN_282 = 8'h19 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_281); // @[FFT.scala 35:12]
  assign _GEN_283 = 8'h1a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_282); // @[FFT.scala 35:12]
  assign _GEN_284 = 8'h1b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_283); // @[FFT.scala 35:12]
  assign _GEN_285 = 8'h1c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_284); // @[FFT.scala 35:12]
  assign _GEN_286 = 8'h1d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_285); // @[FFT.scala 35:12]
  assign _GEN_287 = 8'h1e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_286); // @[FFT.scala 35:12]
  assign _GEN_288 = 8'h1f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_287); // @[FFT.scala 35:12]
  assign _GEN_289 = 8'h20 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_288); // @[FFT.scala 35:12]
  assign _GEN_290 = 8'h21 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_289); // @[FFT.scala 35:12]
  assign _GEN_291 = 8'h22 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_290); // @[FFT.scala 35:12]
  assign _GEN_292 = 8'h23 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_291); // @[FFT.scala 35:12]
  assign _GEN_293 = 8'h24 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_292); // @[FFT.scala 35:12]
  assign _GEN_294 = 8'h25 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_293); // @[FFT.scala 35:12]
  assign _GEN_295 = 8'h26 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_294); // @[FFT.scala 35:12]
  assign _GEN_296 = 8'h27 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_295); // @[FFT.scala 35:12]
  assign _GEN_297 = 8'h28 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_296); // @[FFT.scala 35:12]
  assign _GEN_298 = 8'h29 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_297); // @[FFT.scala 35:12]
  assign _GEN_299 = 8'h2a == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_298); // @[FFT.scala 35:12]
  assign _GEN_300 = 8'h2b == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_299); // @[FFT.scala 35:12]
  assign _GEN_301 = 8'h2c == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_300); // @[FFT.scala 35:12]
  assign _GEN_302 = 8'h2d == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_301); // @[FFT.scala 35:12]
  assign _GEN_303 = 8'h2e == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_302); // @[FFT.scala 35:12]
  assign _GEN_304 = 8'h2f == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_303); // @[FFT.scala 35:12]
  assign _GEN_305 = 8'h30 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_304); // @[FFT.scala 35:12]
  assign _GEN_306 = 8'h31 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_305); // @[FFT.scala 35:12]
  assign _GEN_307 = 8'h32 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_306); // @[FFT.scala 35:12]
  assign _GEN_308 = 8'h33 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_307); // @[FFT.scala 35:12]
  assign _GEN_309 = 8'h34 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_308); // @[FFT.scala 35:12]
  assign _GEN_310 = 8'h35 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_309); // @[FFT.scala 35:12]
  assign _GEN_311 = 8'h36 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_310); // @[FFT.scala 35:12]
  assign _GEN_312 = 8'h37 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_311); // @[FFT.scala 35:12]
  assign _GEN_313 = 8'h38 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_312); // @[FFT.scala 35:12]
  assign _GEN_314 = 8'h39 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_313); // @[FFT.scala 35:12]
  assign _GEN_315 = 8'h3a == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_314); // @[FFT.scala 35:12]
  assign _GEN_316 = 8'h3b == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_315); // @[FFT.scala 35:12]
  assign _GEN_317 = 8'h3c == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_316); // @[FFT.scala 35:12]
  assign _GEN_318 = 8'h3d == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_317); // @[FFT.scala 35:12]
  assign _GEN_319 = 8'h3e == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_318); // @[FFT.scala 35:12]
  assign _GEN_320 = 8'h3f == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_319); // @[FFT.scala 35:12]
  assign _GEN_321 = 8'h40 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_320); // @[FFT.scala 35:12]
  assign _GEN_322 = 8'h41 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_321); // @[FFT.scala 35:12]
  assign _GEN_323 = 8'h42 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_322); // @[FFT.scala 35:12]
  assign _GEN_324 = 8'h43 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_323); // @[FFT.scala 35:12]
  assign _GEN_325 = 8'h44 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_324); // @[FFT.scala 35:12]
  assign _GEN_326 = 8'h45 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_325); // @[FFT.scala 35:12]
  assign _GEN_327 = 8'h46 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_326); // @[FFT.scala 35:12]
  assign _GEN_328 = 8'h47 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_327); // @[FFT.scala 35:12]
  assign _GEN_329 = 8'h48 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_328); // @[FFT.scala 35:12]
  assign _GEN_330 = 8'h49 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_329); // @[FFT.scala 35:12]
  assign _GEN_331 = 8'h4a == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_330); // @[FFT.scala 35:12]
  assign _GEN_332 = 8'h4b == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_331); // @[FFT.scala 35:12]
  assign _GEN_333 = 8'h4c == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_332); // @[FFT.scala 35:12]
  assign _GEN_334 = 8'h4d == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_333); // @[FFT.scala 35:12]
  assign _GEN_335 = 8'h4e == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_334); // @[FFT.scala 35:12]
  assign _GEN_336 = 8'h4f == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_335); // @[FFT.scala 35:12]
  assign _GEN_337 = 8'h50 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_336); // @[FFT.scala 35:12]
  assign _GEN_338 = 8'h51 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_337); // @[FFT.scala 35:12]
  assign _GEN_339 = 8'h52 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_338); // @[FFT.scala 35:12]
  assign _GEN_340 = 8'h53 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_339); // @[FFT.scala 35:12]
  assign _GEN_341 = 8'h54 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_340); // @[FFT.scala 35:12]
  assign _GEN_342 = 8'h55 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_341); // @[FFT.scala 35:12]
  assign _GEN_343 = 8'h56 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_342); // @[FFT.scala 35:12]
  assign _GEN_344 = 8'h57 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_343); // @[FFT.scala 35:12]
  assign _GEN_345 = 8'h58 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_344); // @[FFT.scala 35:12]
  assign _GEN_346 = 8'h59 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_345); // @[FFT.scala 35:12]
  assign _GEN_347 = 8'h5a == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_346); // @[FFT.scala 35:12]
  assign _GEN_348 = 8'h5b == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_347); // @[FFT.scala 35:12]
  assign _GEN_349 = 8'h5c == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_348); // @[FFT.scala 35:12]
  assign _GEN_350 = 8'h5d == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_349); // @[FFT.scala 35:12]
  assign _GEN_351 = 8'h5e == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_350); // @[FFT.scala 35:12]
  assign _GEN_352 = 8'h5f == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_351); // @[FFT.scala 35:12]
  assign _GEN_353 = 8'h60 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_352); // @[FFT.scala 35:12]
  assign _GEN_354 = 8'h61 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_353); // @[FFT.scala 35:12]
  assign _GEN_355 = 8'h62 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_354); // @[FFT.scala 35:12]
  assign _GEN_356 = 8'h63 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_355); // @[FFT.scala 35:12]
  assign _GEN_357 = 8'h64 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_356); // @[FFT.scala 35:12]
  assign _GEN_358 = 8'h65 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_357); // @[FFT.scala 35:12]
  assign _GEN_359 = 8'h66 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_358); // @[FFT.scala 35:12]
  assign _GEN_360 = 8'h67 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_359); // @[FFT.scala 35:12]
  assign _GEN_361 = 8'h68 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_360); // @[FFT.scala 35:12]
  assign _GEN_362 = 8'h69 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_361); // @[FFT.scala 35:12]
  assign _GEN_363 = 8'h6a == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_362); // @[FFT.scala 35:12]
  assign _GEN_364 = 8'h6b == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_363); // @[FFT.scala 35:12]
  assign _GEN_365 = 8'h6c == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_364); // @[FFT.scala 35:12]
  assign _GEN_366 = 8'h6d == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_365); // @[FFT.scala 35:12]
  assign _GEN_367 = 8'h6e == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_366); // @[FFT.scala 35:12]
  assign _GEN_368 = 8'h6f == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_367); // @[FFT.scala 35:12]
  assign _GEN_369 = 8'h70 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_368); // @[FFT.scala 35:12]
  assign _GEN_370 = 8'h71 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_369); // @[FFT.scala 35:12]
  assign _GEN_371 = 8'h72 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_370); // @[FFT.scala 35:12]
  assign _GEN_372 = 8'h73 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_371); // @[FFT.scala 35:12]
  assign _GEN_373 = 8'h74 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_372); // @[FFT.scala 35:12]
  assign _GEN_374 = 8'h75 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_373); // @[FFT.scala 35:12]
  assign _GEN_375 = 8'h76 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_374); // @[FFT.scala 35:12]
  assign _GEN_376 = 8'h77 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_375); // @[FFT.scala 35:12]
  assign _GEN_377 = 8'h78 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_376); // @[FFT.scala 35:12]
  assign _GEN_378 = 8'h79 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_377); // @[FFT.scala 35:12]
  assign _GEN_379 = 8'h7a == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_378); // @[FFT.scala 35:12]
  assign _GEN_380 = 8'h7b == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_379); // @[FFT.scala 35:12]
  assign _GEN_381 = 8'h7c == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_380); // @[FFT.scala 35:12]
  assign _GEN_382 = 8'h7d == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_381); // @[FFT.scala 35:12]
  assign _GEN_383 = 8'h7e == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_382); // @[FFT.scala 35:12]
  assign _GEN_384 = 8'h7f == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_383); // @[FFT.scala 35:12]
  assign _GEN_385 = 8'h80 == cnt[7:0] ? $signed(-32'sh10000) : $signed(_GEN_384); // @[FFT.scala 35:12]
  assign _GEN_386 = 8'h81 == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_385); // @[FFT.scala 35:12]
  assign _GEN_387 = 8'h82 == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_386); // @[FFT.scala 35:12]
  assign _GEN_388 = 8'h83 == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_387); // @[FFT.scala 35:12]
  assign _GEN_389 = 8'h84 == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_388); // @[FFT.scala 35:12]
  assign _GEN_390 = 8'h85 == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_389); // @[FFT.scala 35:12]
  assign _GEN_391 = 8'h86 == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_390); // @[FFT.scala 35:12]
  assign _GEN_392 = 8'h87 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_391); // @[FFT.scala 35:12]
  assign _GEN_393 = 8'h88 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_392); // @[FFT.scala 35:12]
  assign _GEN_394 = 8'h89 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_393); // @[FFT.scala 35:12]
  assign _GEN_395 = 8'h8a == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_394); // @[FFT.scala 35:12]
  assign _GEN_396 = 8'h8b == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_395); // @[FFT.scala 35:12]
  assign _GEN_397 = 8'h8c == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_396); // @[FFT.scala 35:12]
  assign _GEN_398 = 8'h8d == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_397); // @[FFT.scala 35:12]
  assign _GEN_399 = 8'h8e == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_398); // @[FFT.scala 35:12]
  assign _GEN_400 = 8'h8f == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_399); // @[FFT.scala 35:12]
  assign _GEN_401 = 8'h90 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_400); // @[FFT.scala 35:12]
  assign _GEN_402 = 8'h91 == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_401); // @[FFT.scala 35:12]
  assign _GEN_403 = 8'h92 == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_402); // @[FFT.scala 35:12]
  assign _GEN_404 = 8'h93 == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_403); // @[FFT.scala 35:12]
  assign _GEN_405 = 8'h94 == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_404); // @[FFT.scala 35:12]
  assign _GEN_406 = 8'h95 == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_405); // @[FFT.scala 35:12]
  assign _GEN_407 = 8'h96 == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_406); // @[FFT.scala 35:12]
  assign _GEN_408 = 8'h97 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_407); // @[FFT.scala 35:12]
  assign _GEN_409 = 8'h98 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_408); // @[FFT.scala 35:12]
  assign _GEN_410 = 8'h99 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_409); // @[FFT.scala 35:12]
  assign _GEN_411 = 8'h9a == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_410); // @[FFT.scala 35:12]
  assign _GEN_412 = 8'h9b == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_411); // @[FFT.scala 35:12]
  assign _GEN_413 = 8'h9c == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_412); // @[FFT.scala 35:12]
  assign _GEN_414 = 8'h9d == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_413); // @[FFT.scala 35:12]
  assign _GEN_415 = 8'h9e == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_414); // @[FFT.scala 35:12]
  assign _GEN_416 = 8'h9f == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_415); // @[FFT.scala 35:12]
  assign _GEN_417 = 8'ha0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_416); // @[FFT.scala 35:12]
  assign _GEN_418 = 8'ha1 == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_417); // @[FFT.scala 35:12]
  assign _GEN_419 = 8'ha2 == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_418); // @[FFT.scala 35:12]
  assign _GEN_420 = 8'ha3 == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_419); // @[FFT.scala 35:12]
  assign _GEN_421 = 8'ha4 == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_420); // @[FFT.scala 35:12]
  assign _GEN_422 = 8'ha5 == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_421); // @[FFT.scala 35:12]
  assign _GEN_423 = 8'ha6 == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_422); // @[FFT.scala 35:12]
  assign _GEN_424 = 8'ha7 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_423); // @[FFT.scala 35:12]
  assign _GEN_425 = 8'ha8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_424); // @[FFT.scala 35:12]
  assign _GEN_426 = 8'ha9 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_425); // @[FFT.scala 35:12]
  assign _GEN_427 = 8'haa == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_426); // @[FFT.scala 35:12]
  assign _GEN_428 = 8'hab == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_427); // @[FFT.scala 35:12]
  assign _GEN_429 = 8'hac == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_428); // @[FFT.scala 35:12]
  assign _GEN_430 = 8'had == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_429); // @[FFT.scala 35:12]
  assign _GEN_431 = 8'hae == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_430); // @[FFT.scala 35:12]
  assign _GEN_432 = 8'haf == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_431); // @[FFT.scala 35:12]
  assign _GEN_433 = 8'hb0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_432); // @[FFT.scala 35:12]
  assign _GEN_434 = 8'hb1 == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_433); // @[FFT.scala 35:12]
  assign _GEN_435 = 8'hb2 == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_434); // @[FFT.scala 35:12]
  assign _GEN_436 = 8'hb3 == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_435); // @[FFT.scala 35:12]
  assign _GEN_437 = 8'hb4 == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_436); // @[FFT.scala 35:12]
  assign _GEN_438 = 8'hb5 == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_437); // @[FFT.scala 35:12]
  assign _GEN_439 = 8'hb6 == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_438); // @[FFT.scala 35:12]
  assign _GEN_440 = 8'hb7 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_439); // @[FFT.scala 35:12]
  assign _GEN_441 = 8'hb8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_440); // @[FFT.scala 35:12]
  assign _GEN_442 = 8'hb9 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_441); // @[FFT.scala 35:12]
  assign _GEN_443 = 8'hba == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_442); // @[FFT.scala 35:12]
  assign _GEN_444 = 8'hbb == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_443); // @[FFT.scala 35:12]
  assign _GEN_445 = 8'hbc == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_444); // @[FFT.scala 35:12]
  assign _GEN_446 = 8'hbd == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_445); // @[FFT.scala 35:12]
  assign _GEN_447 = 8'hbe == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_446); // @[FFT.scala 35:12]
  assign _GEN_448 = 8'hbf == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_447); // @[FFT.scala 35:12]
  assign _GEN_449 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_448); // @[FFT.scala 35:12]
  assign _GEN_450 = 8'hc1 == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_449); // @[FFT.scala 35:12]
  assign _GEN_451 = 8'hc2 == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_450); // @[FFT.scala 35:12]
  assign _GEN_452 = 8'hc3 == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_451); // @[FFT.scala 35:12]
  assign _GEN_453 = 8'hc4 == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_452); // @[FFT.scala 35:12]
  assign _GEN_454 = 8'hc5 == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_453); // @[FFT.scala 35:12]
  assign _GEN_455 = 8'hc6 == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_454); // @[FFT.scala 35:12]
  assign _GEN_456 = 8'hc7 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_455); // @[FFT.scala 35:12]
  assign _GEN_457 = 8'hc8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_456); // @[FFT.scala 35:12]
  assign _GEN_458 = 8'hc9 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_457); // @[FFT.scala 35:12]
  assign _GEN_459 = 8'hca == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_458); // @[FFT.scala 35:12]
  assign _GEN_460 = 8'hcb == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_459); // @[FFT.scala 35:12]
  assign _GEN_461 = 8'hcc == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_460); // @[FFT.scala 35:12]
  assign _GEN_462 = 8'hcd == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_461); // @[FFT.scala 35:12]
  assign _GEN_463 = 8'hce == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_462); // @[FFT.scala 35:12]
  assign _GEN_464 = 8'hcf == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_463); // @[FFT.scala 35:12]
  assign _GEN_465 = 8'hd0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_464); // @[FFT.scala 35:12]
  assign _GEN_466 = 8'hd1 == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_465); // @[FFT.scala 35:12]
  assign _GEN_467 = 8'hd2 == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_466); // @[FFT.scala 35:12]
  assign _GEN_468 = 8'hd3 == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_467); // @[FFT.scala 35:12]
  assign _GEN_469 = 8'hd4 == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_468); // @[FFT.scala 35:12]
  assign _GEN_470 = 8'hd5 == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_469); // @[FFT.scala 35:12]
  assign _GEN_471 = 8'hd6 == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_470); // @[FFT.scala 35:12]
  assign _GEN_472 = 8'hd7 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_471); // @[FFT.scala 35:12]
  assign _GEN_473 = 8'hd8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_472); // @[FFT.scala 35:12]
  assign _GEN_474 = 8'hd9 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_473); // @[FFT.scala 35:12]
  assign _GEN_475 = 8'hda == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_474); // @[FFT.scala 35:12]
  assign _GEN_476 = 8'hdb == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_475); // @[FFT.scala 35:12]
  assign _GEN_477 = 8'hdc == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_476); // @[FFT.scala 35:12]
  assign _GEN_478 = 8'hdd == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_477); // @[FFT.scala 35:12]
  assign _GEN_479 = 8'hde == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_478); // @[FFT.scala 35:12]
  assign _GEN_480 = 8'hdf == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_479); // @[FFT.scala 35:12]
  assign _GEN_481 = 8'he0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_480); // @[FFT.scala 35:12]
  assign _GEN_482 = 8'he1 == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_481); // @[FFT.scala 35:12]
  assign _GEN_483 = 8'he2 == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_482); // @[FFT.scala 35:12]
  assign _GEN_484 = 8'he3 == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_483); // @[FFT.scala 35:12]
  assign _GEN_485 = 8'he4 == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_484); // @[FFT.scala 35:12]
  assign _GEN_486 = 8'he5 == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_485); // @[FFT.scala 35:12]
  assign _GEN_487 = 8'he6 == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_486); // @[FFT.scala 35:12]
  assign _GEN_488 = 8'he7 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_487); // @[FFT.scala 35:12]
  assign _GEN_489 = 8'he8 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_488); // @[FFT.scala 35:12]
  assign _GEN_490 = 8'he9 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_489); // @[FFT.scala 35:12]
  assign _GEN_491 = 8'hea == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_490); // @[FFT.scala 35:12]
  assign _GEN_492 = 8'heb == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_491); // @[FFT.scala 35:12]
  assign _GEN_493 = 8'hec == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_492); // @[FFT.scala 35:12]
  assign _GEN_494 = 8'hed == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_493); // @[FFT.scala 35:12]
  assign _GEN_495 = 8'hee == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_494); // @[FFT.scala 35:12]
  assign _GEN_496 = 8'hef == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_495); // @[FFT.scala 35:12]
  assign _GEN_497 = 8'hf0 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_496); // @[FFT.scala 35:12]
  assign _GEN_498 = 8'hf1 == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_497); // @[FFT.scala 35:12]
  assign _GEN_499 = 8'hf2 == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_498); // @[FFT.scala 35:12]
  assign _GEN_500 = 8'hf3 == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_499); // @[FFT.scala 35:12]
  assign _GEN_501 = 8'hf4 == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_500); // @[FFT.scala 35:12]
  assign _GEN_502 = 8'hf5 == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_501); // @[FFT.scala 35:12]
  assign _GEN_503 = 8'hf6 == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_502); // @[FFT.scala 35:12]
  assign _GEN_504 = 8'hf7 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_503); // @[FFT.scala 35:12]
  assign _GEN_505 = 8'hf8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_504); // @[FFT.scala 35:12]
  assign _GEN_506 = 8'hf9 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_505); // @[FFT.scala 35:12]
  assign _GEN_507 = 8'hfa == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_506); // @[FFT.scala 35:12]
  assign _GEN_508 = 8'hfb == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_507); // @[FFT.scala 35:12]
  assign _GEN_509 = 8'hfc == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_508); // @[FFT.scala 35:12]
  assign _GEN_510 = 8'hfd == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_509); // @[FFT.scala 35:12]
  assign _GEN_511 = 8'hfe == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_510); // @[FFT.scala 35:12]
  assign _GEN_1282 = 7'h1 == cnt[6:0] ? $signed(32'shffec) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1283 = 7'h2 == cnt[6:0] ? $signed(32'shffb1) : $signed(_GEN_1282); // @[FFT.scala 34:12]
  assign _GEN_1284 = 7'h3 == cnt[6:0] ? $signed(32'shff4e) : $signed(_GEN_1283); // @[FFT.scala 34:12]
  assign _GEN_1285 = 7'h4 == cnt[6:0] ? $signed(32'shfec4) : $signed(_GEN_1284); // @[FFT.scala 34:12]
  assign _GEN_1286 = 7'h5 == cnt[6:0] ? $signed(32'shfe13) : $signed(_GEN_1285); // @[FFT.scala 34:12]
  assign _GEN_1287 = 7'h6 == cnt[6:0] ? $signed(32'shfd3b) : $signed(_GEN_1286); // @[FFT.scala 34:12]
  assign _GEN_1288 = 7'h7 == cnt[6:0] ? $signed(32'shfc3b) : $signed(_GEN_1287); // @[FFT.scala 34:12]
  assign _GEN_1289 = 7'h8 == cnt[6:0] ? $signed(32'shfb15) : $signed(_GEN_1288); // @[FFT.scala 34:12]
  assign _GEN_1290 = 7'h9 == cnt[6:0] ? $signed(32'shf9c8) : $signed(_GEN_1289); // @[FFT.scala 34:12]
  assign _GEN_1291 = 7'ha == cnt[6:0] ? $signed(32'shf854) : $signed(_GEN_1290); // @[FFT.scala 34:12]
  assign _GEN_1292 = 7'hb == cnt[6:0] ? $signed(32'shf6ba) : $signed(_GEN_1291); // @[FFT.scala 34:12]
  assign _GEN_1293 = 7'hc == cnt[6:0] ? $signed(32'shf4fa) : $signed(_GEN_1292); // @[FFT.scala 34:12]
  assign _GEN_1294 = 7'hd == cnt[6:0] ? $signed(32'shf314) : $signed(_GEN_1293); // @[FFT.scala 34:12]
  assign _GEN_1295 = 7'he == cnt[6:0] ? $signed(32'shf109) : $signed(_GEN_1294); // @[FFT.scala 34:12]
  assign _GEN_1296 = 7'hf == cnt[6:0] ? $signed(32'sheed9) : $signed(_GEN_1295); // @[FFT.scala 34:12]
  assign _GEN_1297 = 7'h10 == cnt[6:0] ? $signed(32'shec83) : $signed(_GEN_1296); // @[FFT.scala 34:12]
  assign _GEN_1298 = 7'h11 == cnt[6:0] ? $signed(32'shea0a) : $signed(_GEN_1297); // @[FFT.scala 34:12]
  assign _GEN_1299 = 7'h12 == cnt[6:0] ? $signed(32'she76c) : $signed(_GEN_1298); // @[FFT.scala 34:12]
  assign _GEN_1300 = 7'h13 == cnt[6:0] ? $signed(32'she4aa) : $signed(_GEN_1299); // @[FFT.scala 34:12]
  assign _GEN_1301 = 7'h14 == cnt[6:0] ? $signed(32'she1c6) : $signed(_GEN_1300); // @[FFT.scala 34:12]
  assign _GEN_1302 = 7'h15 == cnt[6:0] ? $signed(32'shdebe) : $signed(_GEN_1301); // @[FFT.scala 34:12]
  assign _GEN_1303 = 7'h16 == cnt[6:0] ? $signed(32'shdb94) : $signed(_GEN_1302); // @[FFT.scala 34:12]
  assign _GEN_1304 = 7'h17 == cnt[6:0] ? $signed(32'shd848) : $signed(_GEN_1303); // @[FFT.scala 34:12]
  assign _GEN_1305 = 7'h18 == cnt[6:0] ? $signed(32'shd4db) : $signed(_GEN_1304); // @[FFT.scala 34:12]
  assign _GEN_1306 = 7'h19 == cnt[6:0] ? $signed(32'shd14d) : $signed(_GEN_1305); // @[FFT.scala 34:12]
  assign _GEN_1307 = 7'h1a == cnt[6:0] ? $signed(32'shcd9f) : $signed(_GEN_1306); // @[FFT.scala 34:12]
  assign _GEN_1308 = 7'h1b == cnt[6:0] ? $signed(32'shc9d1) : $signed(_GEN_1307); // @[FFT.scala 34:12]
  assign _GEN_1309 = 7'h1c == cnt[6:0] ? $signed(32'shc5e4) : $signed(_GEN_1308); // @[FFT.scala 34:12]
  assign _GEN_1310 = 7'h1d == cnt[6:0] ? $signed(32'shc1d8) : $signed(_GEN_1309); // @[FFT.scala 34:12]
  assign _GEN_1311 = 7'h1e == cnt[6:0] ? $signed(32'shbdaf) : $signed(_GEN_1310); // @[FFT.scala 34:12]
  assign _GEN_1312 = 7'h1f == cnt[6:0] ? $signed(32'shb968) : $signed(_GEN_1311); // @[FFT.scala 34:12]
  assign _GEN_1313 = 7'h20 == cnt[6:0] ? $signed(32'shb505) : $signed(_GEN_1312); // @[FFT.scala 34:12]
  assign _GEN_1314 = 7'h21 == cnt[6:0] ? $signed(32'shb086) : $signed(_GEN_1313); // @[FFT.scala 34:12]
  assign _GEN_1315 = 7'h22 == cnt[6:0] ? $signed(32'shabeb) : $signed(_GEN_1314); // @[FFT.scala 34:12]
  assign _GEN_1316 = 7'h23 == cnt[6:0] ? $signed(32'sha736) : $signed(_GEN_1315); // @[FFT.scala 34:12]
  assign _GEN_1317 = 7'h24 == cnt[6:0] ? $signed(32'sha268) : $signed(_GEN_1316); // @[FFT.scala 34:12]
  assign _GEN_1318 = 7'h25 == cnt[6:0] ? $signed(32'sh9d80) : $signed(_GEN_1317); // @[FFT.scala 34:12]
  assign _GEN_1319 = 7'h26 == cnt[6:0] ? $signed(32'sh9880) : $signed(_GEN_1318); // @[FFT.scala 34:12]
  assign _GEN_1320 = 7'h27 == cnt[6:0] ? $signed(32'sh9368) : $signed(_GEN_1319); // @[FFT.scala 34:12]
  assign _GEN_1321 = 7'h28 == cnt[6:0] ? $signed(32'sh8e3a) : $signed(_GEN_1320); // @[FFT.scala 34:12]
  assign _GEN_1322 = 7'h29 == cnt[6:0] ? $signed(32'sh88f6) : $signed(_GEN_1321); // @[FFT.scala 34:12]
  assign _GEN_1323 = 7'h2a == cnt[6:0] ? $signed(32'sh839c) : $signed(_GEN_1322); // @[FFT.scala 34:12]
  assign _GEN_1324 = 7'h2b == cnt[6:0] ? $signed(32'sh7e2f) : $signed(_GEN_1323); // @[FFT.scala 34:12]
  assign _GEN_1325 = 7'h2c == cnt[6:0] ? $signed(32'sh78ad) : $signed(_GEN_1324); // @[FFT.scala 34:12]
  assign _GEN_1326 = 7'h2d == cnt[6:0] ? $signed(32'sh731a) : $signed(_GEN_1325); // @[FFT.scala 34:12]
  assign _GEN_1327 = 7'h2e == cnt[6:0] ? $signed(32'sh6d74) : $signed(_GEN_1326); // @[FFT.scala 34:12]
  assign _GEN_1328 = 7'h2f == cnt[6:0] ? $signed(32'sh67be) : $signed(_GEN_1327); // @[FFT.scala 34:12]
  assign _GEN_1329 = 7'h30 == cnt[6:0] ? $signed(32'sh61f8) : $signed(_GEN_1328); // @[FFT.scala 34:12]
  assign _GEN_1330 = 7'h31 == cnt[6:0] ? $signed(32'sh5c22) : $signed(_GEN_1329); // @[FFT.scala 34:12]
  assign _GEN_1331 = 7'h32 == cnt[6:0] ? $signed(32'sh563e) : $signed(_GEN_1330); // @[FFT.scala 34:12]
  assign _GEN_1332 = 7'h33 == cnt[6:0] ? $signed(32'sh504d) : $signed(_GEN_1331); // @[FFT.scala 34:12]
  assign _GEN_1333 = 7'h34 == cnt[6:0] ? $signed(32'sh4a50) : $signed(_GEN_1332); // @[FFT.scala 34:12]
  assign _GEN_1334 = 7'h35 == cnt[6:0] ? $signed(32'sh4447) : $signed(_GEN_1333); // @[FFT.scala 34:12]
  assign _GEN_1335 = 7'h36 == cnt[6:0] ? $signed(32'sh3e34) : $signed(_GEN_1334); // @[FFT.scala 34:12]
  assign _GEN_1336 = 7'h37 == cnt[6:0] ? $signed(32'sh3817) : $signed(_GEN_1335); // @[FFT.scala 34:12]
  assign _GEN_1337 = 7'h38 == cnt[6:0] ? $signed(32'sh31f1) : $signed(_GEN_1336); // @[FFT.scala 34:12]
  assign _GEN_1338 = 7'h39 == cnt[6:0] ? $signed(32'sh2bc4) : $signed(_GEN_1337); // @[FFT.scala 34:12]
  assign _GEN_1339 = 7'h3a == cnt[6:0] ? $signed(32'sh2590) : $signed(_GEN_1338); // @[FFT.scala 34:12]
  assign _GEN_1340 = 7'h3b == cnt[6:0] ? $signed(32'sh1f56) : $signed(_GEN_1339); // @[FFT.scala 34:12]
  assign _GEN_1341 = 7'h3c == cnt[6:0] ? $signed(32'sh1918) : $signed(_GEN_1340); // @[FFT.scala 34:12]
  assign _GEN_1342 = 7'h3d == cnt[6:0] ? $signed(32'sh12d5) : $signed(_GEN_1341); // @[FFT.scala 34:12]
  assign _GEN_1343 = 7'h3e == cnt[6:0] ? $signed(32'shc90) : $signed(_GEN_1342); // @[FFT.scala 34:12]
  assign _GEN_1344 = 7'h3f == cnt[6:0] ? $signed(32'sh648) : $signed(_GEN_1343); // @[FFT.scala 34:12]
  assign _GEN_1345 = 7'h40 == cnt[6:0] ? $signed(32'sh0) : $signed(_GEN_1344); // @[FFT.scala 34:12]
  assign _GEN_1346 = 7'h41 == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_1345); // @[FFT.scala 34:12]
  assign _GEN_1347 = 7'h42 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_1346); // @[FFT.scala 34:12]
  assign _GEN_1348 = 7'h43 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_1347); // @[FFT.scala 34:12]
  assign _GEN_1349 = 7'h44 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_1348); // @[FFT.scala 34:12]
  assign _GEN_1350 = 7'h45 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_1349); // @[FFT.scala 34:12]
  assign _GEN_1351 = 7'h46 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_1350); // @[FFT.scala 34:12]
  assign _GEN_1352 = 7'h47 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1351); // @[FFT.scala 34:12]
  assign _GEN_1353 = 7'h48 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_1352); // @[FFT.scala 34:12]
  assign _GEN_1354 = 7'h49 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_1353); // @[FFT.scala 34:12]
  assign _GEN_1355 = 7'h4a == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_1354); // @[FFT.scala 34:12]
  assign _GEN_1356 = 7'h4b == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_1355); // @[FFT.scala 34:12]
  assign _GEN_1357 = 7'h4c == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_1356); // @[FFT.scala 34:12]
  assign _GEN_1358 = 7'h4d == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_1357); // @[FFT.scala 34:12]
  assign _GEN_1359 = 7'h4e == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_1358); // @[FFT.scala 34:12]
  assign _GEN_1360 = 7'h4f == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_1359); // @[FFT.scala 34:12]
  assign _GEN_1361 = 7'h50 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_1360); // @[FFT.scala 34:12]
  assign _GEN_1362 = 7'h51 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_1361); // @[FFT.scala 34:12]
  assign _GEN_1363 = 7'h52 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_1362); // @[FFT.scala 34:12]
  assign _GEN_1364 = 7'h53 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_1363); // @[FFT.scala 34:12]
  assign _GEN_1365 = 7'h54 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_1364); // @[FFT.scala 34:12]
  assign _GEN_1366 = 7'h55 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_1365); // @[FFT.scala 34:12]
  assign _GEN_1367 = 7'h56 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_1366); // @[FFT.scala 34:12]
  assign _GEN_1368 = 7'h57 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_1367); // @[FFT.scala 34:12]
  assign _GEN_1369 = 7'h58 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1368); // @[FFT.scala 34:12]
  assign _GEN_1370 = 7'h59 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_1369); // @[FFT.scala 34:12]
  assign _GEN_1371 = 7'h5a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_1370); // @[FFT.scala 34:12]
  assign _GEN_1372 = 7'h5b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_1371); // @[FFT.scala 34:12]
  assign _GEN_1373 = 7'h5c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_1372); // @[FFT.scala 34:12]
  assign _GEN_1374 = 7'h5d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_1373); // @[FFT.scala 34:12]
  assign _GEN_1375 = 7'h5e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_1374); // @[FFT.scala 34:12]
  assign _GEN_1376 = 7'h5f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_1375); // @[FFT.scala 34:12]
  assign _GEN_1377 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_1376); // @[FFT.scala 34:12]
  assign _GEN_1378 = 7'h61 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_1377); // @[FFT.scala 34:12]
  assign _GEN_1379 = 7'h62 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_1378); // @[FFT.scala 34:12]
  assign _GEN_1380 = 7'h63 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_1379); // @[FFT.scala 34:12]
  assign _GEN_1381 = 7'h64 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_1380); // @[FFT.scala 34:12]
  assign _GEN_1382 = 7'h65 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_1381); // @[FFT.scala 34:12]
  assign _GEN_1383 = 7'h66 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_1382); // @[FFT.scala 34:12]
  assign _GEN_1384 = 7'h67 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_1383); // @[FFT.scala 34:12]
  assign _GEN_1385 = 7'h68 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_1384); // @[FFT.scala 34:12]
  assign _GEN_1386 = 7'h69 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_1385); // @[FFT.scala 34:12]
  assign _GEN_1387 = 7'h6a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_1386); // @[FFT.scala 34:12]
  assign _GEN_1388 = 7'h6b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_1387); // @[FFT.scala 34:12]
  assign _GEN_1389 = 7'h6c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_1388); // @[FFT.scala 34:12]
  assign _GEN_1390 = 7'h6d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_1389); // @[FFT.scala 34:12]
  assign _GEN_1391 = 7'h6e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_1390); // @[FFT.scala 34:12]
  assign _GEN_1392 = 7'h6f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_1391); // @[FFT.scala 34:12]
  assign _GEN_1393 = 7'h70 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_1392); // @[FFT.scala 34:12]
  assign _GEN_1394 = 7'h71 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_1393); // @[FFT.scala 34:12]
  assign _GEN_1395 = 7'h72 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_1394); // @[FFT.scala 34:12]
  assign _GEN_1396 = 7'h73 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_1395); // @[FFT.scala 34:12]
  assign _GEN_1397 = 7'h74 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_1396); // @[FFT.scala 34:12]
  assign _GEN_1398 = 7'h75 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_1397); // @[FFT.scala 34:12]
  assign _GEN_1399 = 7'h76 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_1398); // @[FFT.scala 34:12]
  assign _GEN_1400 = 7'h77 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_1399); // @[FFT.scala 34:12]
  assign _GEN_1401 = 7'h78 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_1400); // @[FFT.scala 34:12]
  assign _GEN_1402 = 7'h79 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_1401); // @[FFT.scala 34:12]
  assign _GEN_1403 = 7'h7a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_1402); // @[FFT.scala 34:12]
  assign _GEN_1404 = 7'h7b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_1403); // @[FFT.scala 34:12]
  assign _GEN_1405 = 7'h7c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_1404); // @[FFT.scala 34:12]
  assign _GEN_1406 = 7'h7d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_1405); // @[FFT.scala 34:12]
  assign _GEN_1407 = 7'h7e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_1406); // @[FFT.scala 34:12]
  assign _GEN_1410 = 7'h1 == cnt[6:0] ? $signed(-32'sh648) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1411 = 7'h2 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_1410); // @[FFT.scala 35:12]
  assign _GEN_1412 = 7'h3 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_1411); // @[FFT.scala 35:12]
  assign _GEN_1413 = 7'h4 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_1412); // @[FFT.scala 35:12]
  assign _GEN_1414 = 7'h5 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_1413); // @[FFT.scala 35:12]
  assign _GEN_1415 = 7'h6 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_1414); // @[FFT.scala 35:12]
  assign _GEN_1416 = 7'h7 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1415); // @[FFT.scala 35:12]
  assign _GEN_1417 = 7'h8 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_1416); // @[FFT.scala 35:12]
  assign _GEN_1418 = 7'h9 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_1417); // @[FFT.scala 35:12]
  assign _GEN_1419 = 7'ha == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_1418); // @[FFT.scala 35:12]
  assign _GEN_1420 = 7'hb == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_1419); // @[FFT.scala 35:12]
  assign _GEN_1421 = 7'hc == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_1420); // @[FFT.scala 35:12]
  assign _GEN_1422 = 7'hd == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_1421); // @[FFT.scala 35:12]
  assign _GEN_1423 = 7'he == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_1422); // @[FFT.scala 35:12]
  assign _GEN_1424 = 7'hf == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_1423); // @[FFT.scala 35:12]
  assign _GEN_1425 = 7'h10 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_1424); // @[FFT.scala 35:12]
  assign _GEN_1426 = 7'h11 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_1425); // @[FFT.scala 35:12]
  assign _GEN_1427 = 7'h12 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_1426); // @[FFT.scala 35:12]
  assign _GEN_1428 = 7'h13 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_1427); // @[FFT.scala 35:12]
  assign _GEN_1429 = 7'h14 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_1428); // @[FFT.scala 35:12]
  assign _GEN_1430 = 7'h15 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_1429); // @[FFT.scala 35:12]
  assign _GEN_1431 = 7'h16 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_1430); // @[FFT.scala 35:12]
  assign _GEN_1432 = 7'h17 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_1431); // @[FFT.scala 35:12]
  assign _GEN_1433 = 7'h18 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1432); // @[FFT.scala 35:12]
  assign _GEN_1434 = 7'h19 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_1433); // @[FFT.scala 35:12]
  assign _GEN_1435 = 7'h1a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_1434); // @[FFT.scala 35:12]
  assign _GEN_1436 = 7'h1b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_1435); // @[FFT.scala 35:12]
  assign _GEN_1437 = 7'h1c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_1436); // @[FFT.scala 35:12]
  assign _GEN_1438 = 7'h1d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_1437); // @[FFT.scala 35:12]
  assign _GEN_1439 = 7'h1e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_1438); // @[FFT.scala 35:12]
  assign _GEN_1440 = 7'h1f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_1439); // @[FFT.scala 35:12]
  assign _GEN_1441 = 7'h20 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_1440); // @[FFT.scala 35:12]
  assign _GEN_1442 = 7'h21 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_1441); // @[FFT.scala 35:12]
  assign _GEN_1443 = 7'h22 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_1442); // @[FFT.scala 35:12]
  assign _GEN_1444 = 7'h23 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_1443); // @[FFT.scala 35:12]
  assign _GEN_1445 = 7'h24 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_1444); // @[FFT.scala 35:12]
  assign _GEN_1446 = 7'h25 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_1445); // @[FFT.scala 35:12]
  assign _GEN_1447 = 7'h26 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_1446); // @[FFT.scala 35:12]
  assign _GEN_1448 = 7'h27 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_1447); // @[FFT.scala 35:12]
  assign _GEN_1449 = 7'h28 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_1448); // @[FFT.scala 35:12]
  assign _GEN_1450 = 7'h29 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_1449); // @[FFT.scala 35:12]
  assign _GEN_1451 = 7'h2a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_1450); // @[FFT.scala 35:12]
  assign _GEN_1452 = 7'h2b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_1451); // @[FFT.scala 35:12]
  assign _GEN_1453 = 7'h2c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_1452); // @[FFT.scala 35:12]
  assign _GEN_1454 = 7'h2d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_1453); // @[FFT.scala 35:12]
  assign _GEN_1455 = 7'h2e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_1454); // @[FFT.scala 35:12]
  assign _GEN_1456 = 7'h2f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_1455); // @[FFT.scala 35:12]
  assign _GEN_1457 = 7'h30 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_1456); // @[FFT.scala 35:12]
  assign _GEN_1458 = 7'h31 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_1457); // @[FFT.scala 35:12]
  assign _GEN_1459 = 7'h32 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_1458); // @[FFT.scala 35:12]
  assign _GEN_1460 = 7'h33 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_1459); // @[FFT.scala 35:12]
  assign _GEN_1461 = 7'h34 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_1460); // @[FFT.scala 35:12]
  assign _GEN_1462 = 7'h35 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_1461); // @[FFT.scala 35:12]
  assign _GEN_1463 = 7'h36 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_1462); // @[FFT.scala 35:12]
  assign _GEN_1464 = 7'h37 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_1463); // @[FFT.scala 35:12]
  assign _GEN_1465 = 7'h38 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_1464); // @[FFT.scala 35:12]
  assign _GEN_1466 = 7'h39 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_1465); // @[FFT.scala 35:12]
  assign _GEN_1467 = 7'h3a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_1466); // @[FFT.scala 35:12]
  assign _GEN_1468 = 7'h3b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_1467); // @[FFT.scala 35:12]
  assign _GEN_1469 = 7'h3c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_1468); // @[FFT.scala 35:12]
  assign _GEN_1470 = 7'h3d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_1469); // @[FFT.scala 35:12]
  assign _GEN_1471 = 7'h3e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_1470); // @[FFT.scala 35:12]
  assign _GEN_1472 = 7'h3f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_1471); // @[FFT.scala 35:12]
  assign _GEN_1473 = 7'h40 == cnt[6:0] ? $signed(-32'sh10000) : $signed(_GEN_1472); // @[FFT.scala 35:12]
  assign _GEN_1474 = 7'h41 == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_1473); // @[FFT.scala 35:12]
  assign _GEN_1475 = 7'h42 == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_1474); // @[FFT.scala 35:12]
  assign _GEN_1476 = 7'h43 == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_1475); // @[FFT.scala 35:12]
  assign _GEN_1477 = 7'h44 == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_1476); // @[FFT.scala 35:12]
  assign _GEN_1478 = 7'h45 == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_1477); // @[FFT.scala 35:12]
  assign _GEN_1479 = 7'h46 == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_1478); // @[FFT.scala 35:12]
  assign _GEN_1480 = 7'h47 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_1479); // @[FFT.scala 35:12]
  assign _GEN_1481 = 7'h48 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_1480); // @[FFT.scala 35:12]
  assign _GEN_1482 = 7'h49 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_1481); // @[FFT.scala 35:12]
  assign _GEN_1483 = 7'h4a == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_1482); // @[FFT.scala 35:12]
  assign _GEN_1484 = 7'h4b == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_1483); // @[FFT.scala 35:12]
  assign _GEN_1485 = 7'h4c == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_1484); // @[FFT.scala 35:12]
  assign _GEN_1486 = 7'h4d == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_1485); // @[FFT.scala 35:12]
  assign _GEN_1487 = 7'h4e == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_1486); // @[FFT.scala 35:12]
  assign _GEN_1488 = 7'h4f == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_1487); // @[FFT.scala 35:12]
  assign _GEN_1489 = 7'h50 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_1488); // @[FFT.scala 35:12]
  assign _GEN_1490 = 7'h51 == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_1489); // @[FFT.scala 35:12]
  assign _GEN_1491 = 7'h52 == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_1490); // @[FFT.scala 35:12]
  assign _GEN_1492 = 7'h53 == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_1491); // @[FFT.scala 35:12]
  assign _GEN_1493 = 7'h54 == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_1492); // @[FFT.scala 35:12]
  assign _GEN_1494 = 7'h55 == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_1493); // @[FFT.scala 35:12]
  assign _GEN_1495 = 7'h56 == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_1494); // @[FFT.scala 35:12]
  assign _GEN_1496 = 7'h57 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_1495); // @[FFT.scala 35:12]
  assign _GEN_1497 = 7'h58 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_1496); // @[FFT.scala 35:12]
  assign _GEN_1498 = 7'h59 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_1497); // @[FFT.scala 35:12]
  assign _GEN_1499 = 7'h5a == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_1498); // @[FFT.scala 35:12]
  assign _GEN_1500 = 7'h5b == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_1499); // @[FFT.scala 35:12]
  assign _GEN_1501 = 7'h5c == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_1500); // @[FFT.scala 35:12]
  assign _GEN_1502 = 7'h5d == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_1501); // @[FFT.scala 35:12]
  assign _GEN_1503 = 7'h5e == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_1502); // @[FFT.scala 35:12]
  assign _GEN_1504 = 7'h5f == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_1503); // @[FFT.scala 35:12]
  assign _GEN_1505 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_1504); // @[FFT.scala 35:12]
  assign _GEN_1506 = 7'h61 == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_1505); // @[FFT.scala 35:12]
  assign _GEN_1507 = 7'h62 == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_1506); // @[FFT.scala 35:12]
  assign _GEN_1508 = 7'h63 == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_1507); // @[FFT.scala 35:12]
  assign _GEN_1509 = 7'h64 == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_1508); // @[FFT.scala 35:12]
  assign _GEN_1510 = 7'h65 == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_1509); // @[FFT.scala 35:12]
  assign _GEN_1511 = 7'h66 == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_1510); // @[FFT.scala 35:12]
  assign _GEN_1512 = 7'h67 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_1511); // @[FFT.scala 35:12]
  assign _GEN_1513 = 7'h68 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1512); // @[FFT.scala 35:12]
  assign _GEN_1514 = 7'h69 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_1513); // @[FFT.scala 35:12]
  assign _GEN_1515 = 7'h6a == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_1514); // @[FFT.scala 35:12]
  assign _GEN_1516 = 7'h6b == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_1515); // @[FFT.scala 35:12]
  assign _GEN_1517 = 7'h6c == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_1516); // @[FFT.scala 35:12]
  assign _GEN_1518 = 7'h6d == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_1517); // @[FFT.scala 35:12]
  assign _GEN_1519 = 7'h6e == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_1518); // @[FFT.scala 35:12]
  assign _GEN_1520 = 7'h6f == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_1519); // @[FFT.scala 35:12]
  assign _GEN_1521 = 7'h70 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_1520); // @[FFT.scala 35:12]
  assign _GEN_1522 = 7'h71 == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_1521); // @[FFT.scala 35:12]
  assign _GEN_1523 = 7'h72 == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_1522); // @[FFT.scala 35:12]
  assign _GEN_1524 = 7'h73 == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_1523); // @[FFT.scala 35:12]
  assign _GEN_1525 = 7'h74 == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_1524); // @[FFT.scala 35:12]
  assign _GEN_1526 = 7'h75 == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_1525); // @[FFT.scala 35:12]
  assign _GEN_1527 = 7'h76 == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_1526); // @[FFT.scala 35:12]
  assign _GEN_1528 = 7'h77 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_1527); // @[FFT.scala 35:12]
  assign _GEN_1529 = 7'h78 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_1528); // @[FFT.scala 35:12]
  assign _GEN_1530 = 7'h79 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1529); // @[FFT.scala 35:12]
  assign _GEN_1531 = 7'h7a == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_1530); // @[FFT.scala 35:12]
  assign _GEN_1532 = 7'h7b == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_1531); // @[FFT.scala 35:12]
  assign _GEN_1533 = 7'h7c == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_1532); // @[FFT.scala 35:12]
  assign _GEN_1534 = 7'h7d == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_1533); // @[FFT.scala 35:12]
  assign _GEN_1535 = 7'h7e == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_1534); // @[FFT.scala 35:12]
  assign _GEN_1922 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1923 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_1922); // @[FFT.scala 34:12]
  assign _GEN_1924 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_1923); // @[FFT.scala 34:12]
  assign _GEN_1925 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_1924); // @[FFT.scala 34:12]
  assign _GEN_1926 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_1925); // @[FFT.scala 34:12]
  assign _GEN_1927 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_1926); // @[FFT.scala 34:12]
  assign _GEN_1928 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_1927); // @[FFT.scala 34:12]
  assign _GEN_1929 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_1928); // @[FFT.scala 34:12]
  assign _GEN_1930 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_1929); // @[FFT.scala 34:12]
  assign _GEN_1931 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_1930); // @[FFT.scala 34:12]
  assign _GEN_1932 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_1931); // @[FFT.scala 34:12]
  assign _GEN_1933 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_1932); // @[FFT.scala 34:12]
  assign _GEN_1934 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_1933); // @[FFT.scala 34:12]
  assign _GEN_1935 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_1934); // @[FFT.scala 34:12]
  assign _GEN_1936 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_1935); // @[FFT.scala 34:12]
  assign _GEN_1937 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_1936); // @[FFT.scala 34:12]
  assign _GEN_1938 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_1937); // @[FFT.scala 34:12]
  assign _GEN_1939 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_1938); // @[FFT.scala 34:12]
  assign _GEN_1940 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_1939); // @[FFT.scala 34:12]
  assign _GEN_1941 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_1940); // @[FFT.scala 34:12]
  assign _GEN_1942 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_1941); // @[FFT.scala 34:12]
  assign _GEN_1943 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_1942); // @[FFT.scala 34:12]
  assign _GEN_1944 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_1943); // @[FFT.scala 34:12]
  assign _GEN_1945 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_1944); // @[FFT.scala 34:12]
  assign _GEN_1946 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_1945); // @[FFT.scala 34:12]
  assign _GEN_1947 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_1946); // @[FFT.scala 34:12]
  assign _GEN_1948 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_1947); // @[FFT.scala 34:12]
  assign _GEN_1949 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_1948); // @[FFT.scala 34:12]
  assign _GEN_1950 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_1949); // @[FFT.scala 34:12]
  assign _GEN_1951 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_1950); // @[FFT.scala 34:12]
  assign _GEN_1952 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_1951); // @[FFT.scala 34:12]
  assign _GEN_1953 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_1952); // @[FFT.scala 34:12]
  assign _GEN_1954 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_1953); // @[FFT.scala 34:12]
  assign _GEN_1955 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_1954); // @[FFT.scala 34:12]
  assign _GEN_1956 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_1955); // @[FFT.scala 34:12]
  assign _GEN_1957 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_1956); // @[FFT.scala 34:12]
  assign _GEN_1958 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_1957); // @[FFT.scala 34:12]
  assign _GEN_1959 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_1958); // @[FFT.scala 34:12]
  assign _GEN_1960 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_1959); // @[FFT.scala 34:12]
  assign _GEN_1961 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_1960); // @[FFT.scala 34:12]
  assign _GEN_1962 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_1961); // @[FFT.scala 34:12]
  assign _GEN_1963 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_1962); // @[FFT.scala 34:12]
  assign _GEN_1964 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_1963); // @[FFT.scala 34:12]
  assign _GEN_1965 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1964); // @[FFT.scala 34:12]
  assign _GEN_1966 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_1965); // @[FFT.scala 34:12]
  assign _GEN_1967 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_1966); // @[FFT.scala 34:12]
  assign _GEN_1968 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_1967); // @[FFT.scala 34:12]
  assign _GEN_1969 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_1968); // @[FFT.scala 34:12]
  assign _GEN_1970 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_1969); // @[FFT.scala 34:12]
  assign _GEN_1971 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_1970); // @[FFT.scala 34:12]
  assign _GEN_1972 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_1971); // @[FFT.scala 34:12]
  assign _GEN_1973 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_1972); // @[FFT.scala 34:12]
  assign _GEN_1974 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_1973); // @[FFT.scala 34:12]
  assign _GEN_1975 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_1974); // @[FFT.scala 34:12]
  assign _GEN_1976 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_1975); // @[FFT.scala 34:12]
  assign _GEN_1977 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_1976); // @[FFT.scala 34:12]
  assign _GEN_1978 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_1977); // @[FFT.scala 34:12]
  assign _GEN_1979 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_1978); // @[FFT.scala 34:12]
  assign _GEN_1980 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_1979); // @[FFT.scala 34:12]
  assign _GEN_1981 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_1980); // @[FFT.scala 34:12]
  assign _GEN_1982 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_1981); // @[FFT.scala 34:12]
  assign _GEN_1983 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_1982); // @[FFT.scala 34:12]
  assign _GEN_1986 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1987 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_1986); // @[FFT.scala 35:12]
  assign _GEN_1988 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_1987); // @[FFT.scala 35:12]
  assign _GEN_1989 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_1988); // @[FFT.scala 35:12]
  assign _GEN_1990 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_1989); // @[FFT.scala 35:12]
  assign _GEN_1991 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_1990); // @[FFT.scala 35:12]
  assign _GEN_1992 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_1991); // @[FFT.scala 35:12]
  assign _GEN_1993 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_1992); // @[FFT.scala 35:12]
  assign _GEN_1994 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_1993); // @[FFT.scala 35:12]
  assign _GEN_1995 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_1994); // @[FFT.scala 35:12]
  assign _GEN_1996 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_1995); // @[FFT.scala 35:12]
  assign _GEN_1997 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1996); // @[FFT.scala 35:12]
  assign _GEN_1998 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_1997); // @[FFT.scala 35:12]
  assign _GEN_1999 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_1998); // @[FFT.scala 35:12]
  assign _GEN_2000 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_1999); // @[FFT.scala 35:12]
  assign _GEN_2001 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2000); // @[FFT.scala 35:12]
  assign _GEN_2002 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2001); // @[FFT.scala 35:12]
  assign _GEN_2003 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2002); // @[FFT.scala 35:12]
  assign _GEN_2004 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2003); // @[FFT.scala 35:12]
  assign _GEN_2005 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2004); // @[FFT.scala 35:12]
  assign _GEN_2006 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2005); // @[FFT.scala 35:12]
  assign _GEN_2007 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2006); // @[FFT.scala 35:12]
  assign _GEN_2008 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2007); // @[FFT.scala 35:12]
  assign _GEN_2009 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2008); // @[FFT.scala 35:12]
  assign _GEN_2010 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2009); // @[FFT.scala 35:12]
  assign _GEN_2011 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2010); // @[FFT.scala 35:12]
  assign _GEN_2012 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2011); // @[FFT.scala 35:12]
  assign _GEN_2013 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2012); // @[FFT.scala 35:12]
  assign _GEN_2014 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2013); // @[FFT.scala 35:12]
  assign _GEN_2015 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2014); // @[FFT.scala 35:12]
  assign _GEN_2016 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2015); // @[FFT.scala 35:12]
  assign _GEN_2017 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_2016); // @[FFT.scala 35:12]
  assign _GEN_2018 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2017); // @[FFT.scala 35:12]
  assign _GEN_2019 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2018); // @[FFT.scala 35:12]
  assign _GEN_2020 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2019); // @[FFT.scala 35:12]
  assign _GEN_2021 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2020); // @[FFT.scala 35:12]
  assign _GEN_2022 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2021); // @[FFT.scala 35:12]
  assign _GEN_2023 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2022); // @[FFT.scala 35:12]
  assign _GEN_2024 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2023); // @[FFT.scala 35:12]
  assign _GEN_2025 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2024); // @[FFT.scala 35:12]
  assign _GEN_2026 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2025); // @[FFT.scala 35:12]
  assign _GEN_2027 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2026); // @[FFT.scala 35:12]
  assign _GEN_2028 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2027); // @[FFT.scala 35:12]
  assign _GEN_2029 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2028); // @[FFT.scala 35:12]
  assign _GEN_2030 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2029); // @[FFT.scala 35:12]
  assign _GEN_2031 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2030); // @[FFT.scala 35:12]
  assign _GEN_2032 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2031); // @[FFT.scala 35:12]
  assign _GEN_2033 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2032); // @[FFT.scala 35:12]
  assign _GEN_2034 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2033); // @[FFT.scala 35:12]
  assign _GEN_2035 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2034); // @[FFT.scala 35:12]
  assign _GEN_2036 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2035); // @[FFT.scala 35:12]
  assign _GEN_2037 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2036); // @[FFT.scala 35:12]
  assign _GEN_2038 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2037); // @[FFT.scala 35:12]
  assign _GEN_2039 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2038); // @[FFT.scala 35:12]
  assign _GEN_2040 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2039); // @[FFT.scala 35:12]
  assign _GEN_2041 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2040); // @[FFT.scala 35:12]
  assign _GEN_2042 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2041); // @[FFT.scala 35:12]
  assign _GEN_2043 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2042); // @[FFT.scala 35:12]
  assign _GEN_2044 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2043); // @[FFT.scala 35:12]
  assign _GEN_2045 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2044); // @[FFT.scala 35:12]
  assign _GEN_2046 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2045); // @[FFT.scala 35:12]
  assign _GEN_2047 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2046); // @[FFT.scala 35:12]
  assign _GEN_2242 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_2243 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_2242); // @[FFT.scala 34:12]
  assign _GEN_2244 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_2243); // @[FFT.scala 34:12]
  assign _GEN_2245 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_2244); // @[FFT.scala 34:12]
  assign _GEN_2246 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_2245); // @[FFT.scala 34:12]
  assign _GEN_2247 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_2246); // @[FFT.scala 34:12]
  assign _GEN_2248 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_2247); // @[FFT.scala 34:12]
  assign _GEN_2249 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_2248); // @[FFT.scala 34:12]
  assign _GEN_2250 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_2249); // @[FFT.scala 34:12]
  assign _GEN_2251 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_2250); // @[FFT.scala 34:12]
  assign _GEN_2252 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_2251); // @[FFT.scala 34:12]
  assign _GEN_2253 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_2252); // @[FFT.scala 34:12]
  assign _GEN_2254 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_2253); // @[FFT.scala 34:12]
  assign _GEN_2255 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_2254); // @[FFT.scala 34:12]
  assign _GEN_2256 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_2255); // @[FFT.scala 34:12]
  assign _GEN_2257 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_2256); // @[FFT.scala 34:12]
  assign _GEN_2258 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_2257); // @[FFT.scala 34:12]
  assign _GEN_2259 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_2258); // @[FFT.scala 34:12]
  assign _GEN_2260 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_2259); // @[FFT.scala 34:12]
  assign _GEN_2261 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_2260); // @[FFT.scala 34:12]
  assign _GEN_2262 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_2261); // @[FFT.scala 34:12]
  assign _GEN_2263 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2262); // @[FFT.scala 34:12]
  assign _GEN_2264 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_2263); // @[FFT.scala 34:12]
  assign _GEN_2265 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_2264); // @[FFT.scala 34:12]
  assign _GEN_2266 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_2265); // @[FFT.scala 34:12]
  assign _GEN_2267 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_2266); // @[FFT.scala 34:12]
  assign _GEN_2268 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_2267); // @[FFT.scala 34:12]
  assign _GEN_2269 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_2268); // @[FFT.scala 34:12]
  assign _GEN_2270 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_2269); // @[FFT.scala 34:12]
  assign _GEN_2271 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_2270); // @[FFT.scala 34:12]
  assign _GEN_2274 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_2275 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_2274); // @[FFT.scala 35:12]
  assign _GEN_2276 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_2275); // @[FFT.scala 35:12]
  assign _GEN_2277 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_2276); // @[FFT.scala 35:12]
  assign _GEN_2278 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_2277); // @[FFT.scala 35:12]
  assign _GEN_2279 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2278); // @[FFT.scala 35:12]
  assign _GEN_2280 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_2279); // @[FFT.scala 35:12]
  assign _GEN_2281 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_2280); // @[FFT.scala 35:12]
  assign _GEN_2282 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_2281); // @[FFT.scala 35:12]
  assign _GEN_2283 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_2282); // @[FFT.scala 35:12]
  assign _GEN_2284 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_2283); // @[FFT.scala 35:12]
  assign _GEN_2285 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_2284); // @[FFT.scala 35:12]
  assign _GEN_2286 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_2285); // @[FFT.scala 35:12]
  assign _GEN_2287 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_2286); // @[FFT.scala 35:12]
  assign _GEN_2288 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_2287); // @[FFT.scala 35:12]
  assign _GEN_2289 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_2288); // @[FFT.scala 35:12]
  assign _GEN_2290 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_2289); // @[FFT.scala 35:12]
  assign _GEN_2291 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_2290); // @[FFT.scala 35:12]
  assign _GEN_2292 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_2291); // @[FFT.scala 35:12]
  assign _GEN_2293 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_2292); // @[FFT.scala 35:12]
  assign _GEN_2294 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_2293); // @[FFT.scala 35:12]
  assign _GEN_2295 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_2294); // @[FFT.scala 35:12]
  assign _GEN_2296 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_2295); // @[FFT.scala 35:12]
  assign _GEN_2297 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_2296); // @[FFT.scala 35:12]
  assign _GEN_2298 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_2297); // @[FFT.scala 35:12]
  assign _GEN_2299 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2298); // @[FFT.scala 35:12]
  assign _GEN_2300 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_2299); // @[FFT.scala 35:12]
  assign _GEN_2301 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_2300); // @[FFT.scala 35:12]
  assign _GEN_2302 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_2301); // @[FFT.scala 35:12]
  assign _GEN_2303 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_2302); // @[FFT.scala 35:12]
  assign _GEN_2402 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_2403 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_2402); // @[FFT.scala 34:12]
  assign _GEN_2404 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_2403); // @[FFT.scala 34:12]
  assign _GEN_2405 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_2404); // @[FFT.scala 34:12]
  assign _GEN_2406 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_2405); // @[FFT.scala 34:12]
  assign _GEN_2407 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_2406); // @[FFT.scala 34:12]
  assign _GEN_2408 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_2407); // @[FFT.scala 34:12]
  assign _GEN_2409 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_2408); // @[FFT.scala 34:12]
  assign _GEN_2410 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_2409); // @[FFT.scala 34:12]
  assign _GEN_2411 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_2410); // @[FFT.scala 34:12]
  assign _GEN_2412 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2411); // @[FFT.scala 34:12]
  assign _GEN_2413 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_2412); // @[FFT.scala 34:12]
  assign _GEN_2414 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_2413); // @[FFT.scala 34:12]
  assign _GEN_2415 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_2414); // @[FFT.scala 34:12]
  assign _GEN_2418 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_2419 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_2418); // @[FFT.scala 35:12]
  assign _GEN_2420 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2419); // @[FFT.scala 35:12]
  assign _GEN_2421 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_2420); // @[FFT.scala 35:12]
  assign _GEN_2422 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_2421); // @[FFT.scala 35:12]
  assign _GEN_2423 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_2422); // @[FFT.scala 35:12]
  assign _GEN_2424 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_2423); // @[FFT.scala 35:12]
  assign _GEN_2425 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_2424); // @[FFT.scala 35:12]
  assign _GEN_2426 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_2425); // @[FFT.scala 35:12]
  assign _GEN_2427 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_2426); // @[FFT.scala 35:12]
  assign _GEN_2428 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_2427); // @[FFT.scala 35:12]
  assign _GEN_2429 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_2428); // @[FFT.scala 35:12]
  assign _GEN_2430 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2429); // @[FFT.scala 35:12]
  assign _GEN_2431 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_2430); // @[FFT.scala 35:12]
  assign _GEN_2482 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_2483 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_2482); // @[FFT.scala 34:12]
  assign _GEN_2484 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_2483); // @[FFT.scala 34:12]
  assign _GEN_2485 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_2484); // @[FFT.scala 34:12]
  assign _GEN_2486 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_2485); // @[FFT.scala 34:12]
  assign _GEN_2487 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_2486); // @[FFT.scala 34:12]
  assign _GEN_2490 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_2491 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_2490); // @[FFT.scala 35:12]
  assign _GEN_2492 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_2491); // @[FFT.scala 35:12]
  assign _GEN_2493 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_2492); // @[FFT.scala 35:12]
  assign _GEN_2494 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_2493); // @[FFT.scala 35:12]
  assign _GEN_2495 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_2494); // @[FFT.scala 35:12]
  assign _GEN_2522 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_2523 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_2522); // @[FFT.scala 34:12]
  assign _GEN_2526 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_2527 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_2526); // @[FFT.scala 35:12]
  assign io_dOut1_re = _T_947_re; // @[FFT.scala 62:12]
  assign io_dOut1_im = _T_947_im; // @[FFT.scala 62:12]
  assign io_dOut2_re = _T_948_re; // @[FFT.scala 63:12]
  assign io_dOut2_im = _T_948_im; // @[FFT.scala 63:12]
  assign io_dout_valid = _T_1460; // @[FFT.scala 64:17]
  assign Butterfly_io_in1_re = _T_401_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_401_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = io_dIn_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = 8'hff == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_255); // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = 8'hff == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_511); // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_530_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_530_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cnt[7]; // @[Butterfly.scala 113:17]
  assign Butterfly_1_io_in1_re = _T_662_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_662_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = 7'h7f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_1407); // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = 7'h7f == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_1535); // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_727_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_727_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cnt[6]; // @[Butterfly.scala 113:17]
  assign Butterfly_2_io_in1_re = _T_795_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_795_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_1983); // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_2047); // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_828_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_828_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cnt[5]; // @[Butterfly.scala 113:17]
  assign Butterfly_3_io_in1_re = _T_864_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_864_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_2271); // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_2303); // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_881_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_881_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cnt[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_901_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_901_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_2415); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_2431); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_910_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_910_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cnt[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_922_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_922_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_2487); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_2495); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_927_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_927_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cnt[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_935_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_935_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_2523); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_2527); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_938_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_938_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cnt[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_7_io_in1_re = _T_944_re; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in1_im = _T_944_im; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_7_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in2_re = _T_946_re; // @[Butterfly.scala 112:17]
  assign Switch_7_io_in2_im = _T_946_im; // @[Butterfly.scala 112:17]
  assign Switch_7_io_sel = cnt[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_146_re = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146_im = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_147_re = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_147_im = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_148_re = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_148_im = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_149_re = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_149_im = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_150_re = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_150_im = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_151_re = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_151_im = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_152_re = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_152_im = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_153_re = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_153_im = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_154_re = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_154_im = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_155_re = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_155_im = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_156_re = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_156_im = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_157_re = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_157_im = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_158_re = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_158_im = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_159_re = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_159_im = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_160_re = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_160_im = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_161_re = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_161_im = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_162_re = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_162_im = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_163_re = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_163_im = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_164_re = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_164_im = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_165_re = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_165_im = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_166_re = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_166_im = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_167_re = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_167_im = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_168_re = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_168_im = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_169_re = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_169_im = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_170_re = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_170_im = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_171_re = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_171_im = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_172_re = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_172_im = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_173_re = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_173_im = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_174_re = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_174_im = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_175_re = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_175_im = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_176_re = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_176_im = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_177_re = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_177_im = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_178_re = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_178_im = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_179_re = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_179_im = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_180_re = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_180_im = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_181_re = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_181_im = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_182_re = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_182_im = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_183_re = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_183_im = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_184_re = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_184_im = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_185_re = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_185_im = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_186_re = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_186_im = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_187_re = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_187_im = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_188_re = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_188_im = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_189_re = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_189_im = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_190_re = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_190_im = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_191_re = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_191_im = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_192_re = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_192_im = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_193_re = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_193_im = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_194_re = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_194_im = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_195_re = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_195_im = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_196_re = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_196_im = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_197_re = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_197_im = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_198_re = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_198_im = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_199_re = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_199_im = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_200_re = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_200_im = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_201_re = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_201_im = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_202_re = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_202_im = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_203_re = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_203_im = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_204_re = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_204_im = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_205_re = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_205_im = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_206_re = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_206_im = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_207_re = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_207_im = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_208_re = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_208_im = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_209_re = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_209_im = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_210_re = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_210_im = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_211_re = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_211_im = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_212_re = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_212_im = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_213_re = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_213_im = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_214_re = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_214_im = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_215_re = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_215_im = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_216_re = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_216_im = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_217_re = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_217_im = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_218_re = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_218_im = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_219_re = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_219_im = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_220_re = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_220_im = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_221_re = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_221_im = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_222_re = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_222_im = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_223_re = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_223_im = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_224_re = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_224_im = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_225_re = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_225_im = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_226_re = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_226_im = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_227_re = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_227_im = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_228_re = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_228_im = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_229_re = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_229_im = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_230_re = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_230_im = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_231_re = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_231_im = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_232_re = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_232_im = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_233_re = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_233_im = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_234_re = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_234_im = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_235_re = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_235_im = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_236_re = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_236_im = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_237_re = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_237_im = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_238_re = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_238_im = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_239_re = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_239_im = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_240_re = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_240_im = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_241_re = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_241_im = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_242_re = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_242_im = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_243_re = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_243_im = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_244_re = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_244_im = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_245_re = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_245_im = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_246_re = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_246_im = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_247_re = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_247_im = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_248_re = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_248_im = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_249_re = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_249_im = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_250_re = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_250_im = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_251_re = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_251_im = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_252_re = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_252_im = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_253_re = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_253_im = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_254_re = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_254_im = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_255_re = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_255_im = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_256_re = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_256_im = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_257_re = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_257_im = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_258_re = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_258_im = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_259_re = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_259_im = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_260_re = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_260_im = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_261_re = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_261_im = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_262_re = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_262_im = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_263_re = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_263_im = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_264_re = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_264_im = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_265_re = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_265_im = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_266_re = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_266_im = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_267_re = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_267_im = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_268_re = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_268_im = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_269_re = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_269_im = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_270_re = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_270_im = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_271_re = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_271_im = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_272_re = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_272_im = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_273_re = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_273_im = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_274_re = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_274_im = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_275_re = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_275_im = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_276_re = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_276_im = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_277_re = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_277_im = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_278_re = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_278_im = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_279_re = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_279_im = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_280_re = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_280_im = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_281_re = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_281_im = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_282_re = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_282_im = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_283_re = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_283_im = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_284_re = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_284_im = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_285_re = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_285_im = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_286_re = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_286_im = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_287_re = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_287_im = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_288_re = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_288_im = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_289_re = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_289_im = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_290_re = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_290_im = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_291_re = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_291_im = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_292_re = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_292_im = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_293_re = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_293_im = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_294_re = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_294_im = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_295_re = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_295_im = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_296_re = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_296_im = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_297_re = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_297_im = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_298_re = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_298_im = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_299_re = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_299_im = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_300_re = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_300_im = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_301_re = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_301_im = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_302_re = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_302_im = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_303_re = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_303_im = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_304_re = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_304_im = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_305_re = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_305_im = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_306_re = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_306_im = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_307_re = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_307_im = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_308_re = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_308_im = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_309_re = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_309_im = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_310_re = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_310_im = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_311_re = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_311_im = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_312_re = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_312_im = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_313_re = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_313_im = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_314_re = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_314_im = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_315_re = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_315_im = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_316_re = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_316_im = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_317_re = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_317_im = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_318_re = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_318_im = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_319_re = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_319_im = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_320_re = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_320_im = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_321_re = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_321_im = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_322_re = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_322_im = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_323_re = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_323_im = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_324_re = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_324_im = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_325_re = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_325_im = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_326_re = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_326_im = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_327_re = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_327_im = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_328_re = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_328_im = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_329_re = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_329_im = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_330_re = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_330_im = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_331_re = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_331_im = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_332_re = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_332_im = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_333_re = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_333_im = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_334_re = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_334_im = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_335_re = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_335_im = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_336_re = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_336_im = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_337_re = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_337_im = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_338_re = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_338_im = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_339_re = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_339_im = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_340_re = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_340_im = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_341_re = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_341_im = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_342_re = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_342_im = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_343_re = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_343_im = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_344_re = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_344_im = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_345_re = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_345_im = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_346_re = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_346_im = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_347_re = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_347_im = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_348_re = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_348_im = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_349_re = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_349_im = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_350_re = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_350_im = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_351_re = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_351_im = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_352_re = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_352_im = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_353_re = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_353_im = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_354_re = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_354_im = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_355_re = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_355_im = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_356_re = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_356_im = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_357_re = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_357_im = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_358_re = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_358_im = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_359_re = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_359_im = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_360_re = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_360_im = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_361_re = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_361_im = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_362_re = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_362_im = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_363_re = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_363_im = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_364_re = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_364_im = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_365_re = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_365_im = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_366_re = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_366_im = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_367_re = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_367_im = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_368_re = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_368_im = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_369_re = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_369_im = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_370_re = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_370_im = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_371_re = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_371_im = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_372_re = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_372_im = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_373_re = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_373_im = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_374_re = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_374_im = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_375_re = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_375_im = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_376_re = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_376_im = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_377_re = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_377_im = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_378_re = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_378_im = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_379_re = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_379_im = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_380_re = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_380_im = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_381_re = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_381_im = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_382_re = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_382_im = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_383_re = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_383_im = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_384_re = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_384_im = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_385_re = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_385_im = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_386_re = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_386_im = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_387_re = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_387_im = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_388_re = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_388_im = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_389_re = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_389_im = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_390_re = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_390_im = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_391_re = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_391_im = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_392_re = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_392_im = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_393_re = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_393_im = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_394_re = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_394_im = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_395_re = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_395_im = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_396_re = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_396_im = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_397_re = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_397_im = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_398_re = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_398_im = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_399_re = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_399_im = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_400_re = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_400_im = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_401_re = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_401_im = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_403_re = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_403_im = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_404_re = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_404_im = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_405_re = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_405_im = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_406_re = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_406_im = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_407_re = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_407_im = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_408_re = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_408_im = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_409_re = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_409_im = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_410_re = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_410_im = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_411_re = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_411_im = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_412_re = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_412_im = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_413_re = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_413_im = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_414_re = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_414_im = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_415_re = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_415_im = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_416_re = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_416_im = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_417_re = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_417_im = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_418_re = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_418_im = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_419_re = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_419_im = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_420_re = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_420_im = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_421_re = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_421_im = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_422_re = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_422_im = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_423_re = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_423_im = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_424_re = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_424_im = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_425_re = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_425_im = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_426_re = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_426_im = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_427_re = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_427_im = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_428_re = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_428_im = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_429_re = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_429_im = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_430_re = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_430_im = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_431_re = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_431_im = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_432_re = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_432_im = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_433_re = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_433_im = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_434_re = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_434_im = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_435_re = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_435_im = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_436_re = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_436_im = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_437_re = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_437_im = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_438_re = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_438_im = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_439_re = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_439_im = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_440_re = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_440_im = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_441_re = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_441_im = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_442_re = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_442_im = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_443_re = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_443_im = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_444_re = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_444_im = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_445_re = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_445_im = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_446_re = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_446_im = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_447_re = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_447_im = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_448_re = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_448_im = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_449_re = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_449_im = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_450_re = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_450_im = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_451_re = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_451_im = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_452_re = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_452_im = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_453_re = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_453_im = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_454_re = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_454_im = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_455_re = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_455_im = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_456_re = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_456_im = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_457_re = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_457_im = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_458_re = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_458_im = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_459_re = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_459_im = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_460_re = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_460_im = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_461_re = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_461_im = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_462_re = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_462_im = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_463_re = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_463_im = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_464_re = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_464_im = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_465_re = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_465_im = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_466_re = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_466_im = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_467_re = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_467_im = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_468_re = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_468_im = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_469_re = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_469_im = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_470_re = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_470_im = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_471_re = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_471_im = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_472_re = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_472_im = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_473_re = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_473_im = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_474_re = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_474_im = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_475_re = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_475_im = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_476_re = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_476_im = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_477_re = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_477_im = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_478_re = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_478_im = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_479_re = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_479_im = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_480_re = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_480_im = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_481_re = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_481_im = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_482_re = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_482_im = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_483_re = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_483_im = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_484_re = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_484_im = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_485_re = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_485_im = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_486_re = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_486_im = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_487_re = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_487_im = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_488_re = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_488_im = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_489_re = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_489_im = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_490_re = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_490_im = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_491_re = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_491_im = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_492_re = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_492_im = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_493_re = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_493_im = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_494_re = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_494_im = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_495_re = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_495_im = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_496_re = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_496_im = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_497_re = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_497_im = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_498_re = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_498_im = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_499_re = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_499_im = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_500_re = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_500_im = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_501_re = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_501_im = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_502_re = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_502_im = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_503_re = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_503_im = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_504_re = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_504_im = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_505_re = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_505_im = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_506_re = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_506_im = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_507_re = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_507_im = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_508_re = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_508_im = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_509_re = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_509_im = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_510_re = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_510_im = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_511_re = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_511_im = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_512_re = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_512_im = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_513_re = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_513_im = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_514_re = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_514_im = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_515_re = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_515_im = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_516_re = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_516_im = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_517_re = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_517_im = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_518_re = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_518_im = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_519_re = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_519_im = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_520_re = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_520_im = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_521_re = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_521_im = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_522_re = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_522_im = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_523_re = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_523_im = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_524_re = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_524_im = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_525_re = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_525_im = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_526_re = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_526_im = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_527_re = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_527_im = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_528_re = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_528_im = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_529_re = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_529_im = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_530_re = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_530_im = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_535_re = _RAND_769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_535_im = _RAND_770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_536_re = _RAND_771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_536_im = _RAND_772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_537_re = _RAND_773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_537_im = _RAND_774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_538_re = _RAND_775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_538_im = _RAND_776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_539_re = _RAND_777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_539_im = _RAND_778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_540_re = _RAND_779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_540_im = _RAND_780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_541_re = _RAND_781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_541_im = _RAND_782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_542_re = _RAND_783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_542_im = _RAND_784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_543_re = _RAND_785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_543_im = _RAND_786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_544_re = _RAND_787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_544_im = _RAND_788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_545_re = _RAND_789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_545_im = _RAND_790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_546_re = _RAND_791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_546_im = _RAND_792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_547_re = _RAND_793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_547_im = _RAND_794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_548_re = _RAND_795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_548_im = _RAND_796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_549_re = _RAND_797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_549_im = _RAND_798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_550_re = _RAND_799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_550_im = _RAND_800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_551_re = _RAND_801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_551_im = _RAND_802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_552_re = _RAND_803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_552_im = _RAND_804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_553_re = _RAND_805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_553_im = _RAND_806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_554_re = _RAND_807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_554_im = _RAND_808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_555_re = _RAND_809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_555_im = _RAND_810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_556_re = _RAND_811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_556_im = _RAND_812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_557_re = _RAND_813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_557_im = _RAND_814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_558_re = _RAND_815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_558_im = _RAND_816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_559_re = _RAND_817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_559_im = _RAND_818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_560_re = _RAND_819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_560_im = _RAND_820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_561_re = _RAND_821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_561_im = _RAND_822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_562_re = _RAND_823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_562_im = _RAND_824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_563_re = _RAND_825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_563_im = _RAND_826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_564_re = _RAND_827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_564_im = _RAND_828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_565_re = _RAND_829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_565_im = _RAND_830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_566_re = _RAND_831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_566_im = _RAND_832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_567_re = _RAND_833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_567_im = _RAND_834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_568_re = _RAND_835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_568_im = _RAND_836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_569_re = _RAND_837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_569_im = _RAND_838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_570_re = _RAND_839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_570_im = _RAND_840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_571_re = _RAND_841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_571_im = _RAND_842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_572_re = _RAND_843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_572_im = _RAND_844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_573_re = _RAND_845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_573_im = _RAND_846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_574_re = _RAND_847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_574_im = _RAND_848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_575_re = _RAND_849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_575_im = _RAND_850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_576_re = _RAND_851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_576_im = _RAND_852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_577_re = _RAND_853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_577_im = _RAND_854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_578_re = _RAND_855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_578_im = _RAND_856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_579_re = _RAND_857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_579_im = _RAND_858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_580_re = _RAND_859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_580_im = _RAND_860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_581_re = _RAND_861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_581_im = _RAND_862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_582_re = _RAND_863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_582_im = _RAND_864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_583_re = _RAND_865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_583_im = _RAND_866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_584_re = _RAND_867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_584_im = _RAND_868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_585_re = _RAND_869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_585_im = _RAND_870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_586_re = _RAND_871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_586_im = _RAND_872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_587_re = _RAND_873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_587_im = _RAND_874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_588_re = _RAND_875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_588_im = _RAND_876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_589_re = _RAND_877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_589_im = _RAND_878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_590_re = _RAND_879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_590_im = _RAND_880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_591_re = _RAND_881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_591_im = _RAND_882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_592_re = _RAND_883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_592_im = _RAND_884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_593_re = _RAND_885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_593_im = _RAND_886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_594_re = _RAND_887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_594_im = _RAND_888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_595_re = _RAND_889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_595_im = _RAND_890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_596_re = _RAND_891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_596_im = _RAND_892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_597_re = _RAND_893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_597_im = _RAND_894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_598_re = _RAND_895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_598_im = _RAND_896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_599_re = _RAND_897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_599_im = _RAND_898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_600_re = _RAND_899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_600_im = _RAND_900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_601_re = _RAND_901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_601_im = _RAND_902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_602_re = _RAND_903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_602_im = _RAND_904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_603_re = _RAND_905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_603_im = _RAND_906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_604_re = _RAND_907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_604_im = _RAND_908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_605_re = _RAND_909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_605_im = _RAND_910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_606_re = _RAND_911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_606_im = _RAND_912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_607_re = _RAND_913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_607_im = _RAND_914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_608_re = _RAND_915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_608_im = _RAND_916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_609_re = _RAND_917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_609_im = _RAND_918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_610_re = _RAND_919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_610_im = _RAND_920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_611_re = _RAND_921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_611_im = _RAND_922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_612_re = _RAND_923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_612_im = _RAND_924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_613_re = _RAND_925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_613_im = _RAND_926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_614_re = _RAND_927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_614_im = _RAND_928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_615_re = _RAND_929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_615_im = _RAND_930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_616_re = _RAND_931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_616_im = _RAND_932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_617_re = _RAND_933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_617_im = _RAND_934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_618_re = _RAND_935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_618_im = _RAND_936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_619_re = _RAND_937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_619_im = _RAND_938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_620_re = _RAND_939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_620_im = _RAND_940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_621_re = _RAND_941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_621_im = _RAND_942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_622_re = _RAND_943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_622_im = _RAND_944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_623_re = _RAND_945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_623_im = _RAND_946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_624_re = _RAND_947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_624_im = _RAND_948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_625_re = _RAND_949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_625_im = _RAND_950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_626_re = _RAND_951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_626_im = _RAND_952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_627_re = _RAND_953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_627_im = _RAND_954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_628_re = _RAND_955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_628_im = _RAND_956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_629_re = _RAND_957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_629_im = _RAND_958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_630_re = _RAND_959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_630_im = _RAND_960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_631_re = _RAND_961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_631_im = _RAND_962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_632_re = _RAND_963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_632_im = _RAND_964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_633_re = _RAND_965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_633_im = _RAND_966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_634_re = _RAND_967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_634_im = _RAND_968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_635_re = _RAND_969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_635_im = _RAND_970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_636_re = _RAND_971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_636_im = _RAND_972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_637_re = _RAND_973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_637_im = _RAND_974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_638_re = _RAND_975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_638_im = _RAND_976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_639_re = _RAND_977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_639_im = _RAND_978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_640_re = _RAND_979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_640_im = _RAND_980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_641_re = _RAND_981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_641_im = _RAND_982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_642_re = _RAND_983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_642_im = _RAND_984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_643_re = _RAND_985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_643_im = _RAND_986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_644_re = _RAND_987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_644_im = _RAND_988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_645_re = _RAND_989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_645_im = _RAND_990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_646_re = _RAND_991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_646_im = _RAND_992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_647_re = _RAND_993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_647_im = _RAND_994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_648_re = _RAND_995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_648_im = _RAND_996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_649_re = _RAND_997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_649_im = _RAND_998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_650_re = _RAND_999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_650_im = _RAND_1000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_651_re = _RAND_1001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_651_im = _RAND_1002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_652_re = _RAND_1003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_652_im = _RAND_1004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_653_re = _RAND_1005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_653_im = _RAND_1006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_654_re = _RAND_1007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_654_im = _RAND_1008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_655_re = _RAND_1009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_655_im = _RAND_1010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_656_re = _RAND_1011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_656_im = _RAND_1012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_657_re = _RAND_1013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_657_im = _RAND_1014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_658_re = _RAND_1015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_658_im = _RAND_1016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_659_re = _RAND_1017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_659_im = _RAND_1018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_660_re = _RAND_1019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_660_im = _RAND_1020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_661_re = _RAND_1021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_661_im = _RAND_1022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_662_re = _RAND_1023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_662_im = _RAND_1024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_664_re = _RAND_1025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_664_im = _RAND_1026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_665_re = _RAND_1027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_665_im = _RAND_1028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_666_re = _RAND_1029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_666_im = _RAND_1030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_667_re = _RAND_1031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_667_im = _RAND_1032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_668_re = _RAND_1033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_668_im = _RAND_1034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_669_re = _RAND_1035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_669_im = _RAND_1036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_670_re = _RAND_1037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_670_im = _RAND_1038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_671_re = _RAND_1039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_671_im = _RAND_1040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_672_re = _RAND_1041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_672_im = _RAND_1042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_673_re = _RAND_1043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_673_im = _RAND_1044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_674_re = _RAND_1045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_674_im = _RAND_1046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_675_re = _RAND_1047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_675_im = _RAND_1048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_676_re = _RAND_1049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_676_im = _RAND_1050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_677_re = _RAND_1051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_677_im = _RAND_1052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_678_re = _RAND_1053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_678_im = _RAND_1054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_679_re = _RAND_1055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_679_im = _RAND_1056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_680_re = _RAND_1057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_680_im = _RAND_1058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_681_re = _RAND_1059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_681_im = _RAND_1060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_682_re = _RAND_1061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_682_im = _RAND_1062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_683_re = _RAND_1063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_683_im = _RAND_1064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_684_re = _RAND_1065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_684_im = _RAND_1066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_685_re = _RAND_1067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_685_im = _RAND_1068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_686_re = _RAND_1069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_686_im = _RAND_1070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_687_re = _RAND_1071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_687_im = _RAND_1072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_688_re = _RAND_1073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_688_im = _RAND_1074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_689_re = _RAND_1075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_689_im = _RAND_1076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_690_re = _RAND_1077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_690_im = _RAND_1078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_691_re = _RAND_1079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_691_im = _RAND_1080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_692_re = _RAND_1081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_692_im = _RAND_1082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_693_re = _RAND_1083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_693_im = _RAND_1084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_694_re = _RAND_1085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_694_im = _RAND_1086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_695_re = _RAND_1087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_695_im = _RAND_1088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_696_re = _RAND_1089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_696_im = _RAND_1090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_697_re = _RAND_1091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_697_im = _RAND_1092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_698_re = _RAND_1093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_698_im = _RAND_1094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_699_re = _RAND_1095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_699_im = _RAND_1096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_700_re = _RAND_1097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_700_im = _RAND_1098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_701_re = _RAND_1099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_701_im = _RAND_1100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_702_re = _RAND_1101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_702_im = _RAND_1102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_703_re = _RAND_1103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_703_im = _RAND_1104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_704_re = _RAND_1105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_704_im = _RAND_1106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_705_re = _RAND_1107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_705_im = _RAND_1108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_706_re = _RAND_1109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_706_im = _RAND_1110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_707_re = _RAND_1111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_707_im = _RAND_1112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_708_re = _RAND_1113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_708_im = _RAND_1114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_709_re = _RAND_1115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_709_im = _RAND_1116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_710_re = _RAND_1117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_710_im = _RAND_1118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_711_re = _RAND_1119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_711_im = _RAND_1120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_712_re = _RAND_1121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_712_im = _RAND_1122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_713_re = _RAND_1123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_713_im = _RAND_1124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_714_re = _RAND_1125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_714_im = _RAND_1126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_715_re = _RAND_1127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_715_im = _RAND_1128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_716_re = _RAND_1129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_716_im = _RAND_1130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_717_re = _RAND_1131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_717_im = _RAND_1132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_718_re = _RAND_1133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_718_im = _RAND_1134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_719_re = _RAND_1135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_719_im = _RAND_1136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_720_re = _RAND_1137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_720_im = _RAND_1138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_721_re = _RAND_1139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_721_im = _RAND_1140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_722_re = _RAND_1141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_722_im = _RAND_1142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_723_re = _RAND_1143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_723_im = _RAND_1144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_724_re = _RAND_1145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_724_im = _RAND_1146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_725_re = _RAND_1147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_725_im = _RAND_1148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_726_re = _RAND_1149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_726_im = _RAND_1150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_727_re = _RAND_1151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_727_im = _RAND_1152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_732_re = _RAND_1153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_732_im = _RAND_1154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_733_re = _RAND_1155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_733_im = _RAND_1156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_734_re = _RAND_1157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_734_im = _RAND_1158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_735_re = _RAND_1159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_735_im = _RAND_1160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_736_re = _RAND_1161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_736_im = _RAND_1162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_737_re = _RAND_1163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_737_im = _RAND_1164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_738_re = _RAND_1165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_738_im = _RAND_1166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_739_re = _RAND_1167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_739_im = _RAND_1168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_740_re = _RAND_1169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_740_im = _RAND_1170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_741_re = _RAND_1171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_741_im = _RAND_1172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_742_re = _RAND_1173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_742_im = _RAND_1174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_743_re = _RAND_1175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_743_im = _RAND_1176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_744_re = _RAND_1177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_744_im = _RAND_1178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_745_re = _RAND_1179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_745_im = _RAND_1180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_746_re = _RAND_1181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_746_im = _RAND_1182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_747_re = _RAND_1183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_747_im = _RAND_1184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_748_re = _RAND_1185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_748_im = _RAND_1186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_749_re = _RAND_1187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_749_im = _RAND_1188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_750_re = _RAND_1189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_750_im = _RAND_1190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_751_re = _RAND_1191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_751_im = _RAND_1192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_752_re = _RAND_1193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_752_im = _RAND_1194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_753_re = _RAND_1195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_753_im = _RAND_1196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_754_re = _RAND_1197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_754_im = _RAND_1198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_755_re = _RAND_1199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_755_im = _RAND_1200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_756_re = _RAND_1201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_756_im = _RAND_1202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_757_re = _RAND_1203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_757_im = _RAND_1204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_758_re = _RAND_1205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_758_im = _RAND_1206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_759_re = _RAND_1207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_759_im = _RAND_1208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_760_re = _RAND_1209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_760_im = _RAND_1210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_761_re = _RAND_1211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_761_im = _RAND_1212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_762_re = _RAND_1213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_762_im = _RAND_1214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_763_re = _RAND_1215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_763_im = _RAND_1216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_764_re = _RAND_1217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_764_im = _RAND_1218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_765_re = _RAND_1219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_765_im = _RAND_1220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_766_re = _RAND_1221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_766_im = _RAND_1222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_767_re = _RAND_1223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_767_im = _RAND_1224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_768_re = _RAND_1225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_768_im = _RAND_1226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_769_re = _RAND_1227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_769_im = _RAND_1228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_770_re = _RAND_1229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_770_im = _RAND_1230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_771_re = _RAND_1231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_771_im = _RAND_1232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_772_re = _RAND_1233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_772_im = _RAND_1234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_773_re = _RAND_1235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_773_im = _RAND_1236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_774_re = _RAND_1237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_774_im = _RAND_1238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_775_re = _RAND_1239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_775_im = _RAND_1240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_776_re = _RAND_1241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_776_im = _RAND_1242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_777_re = _RAND_1243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_777_im = _RAND_1244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_778_re = _RAND_1245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_778_im = _RAND_1246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_779_re = _RAND_1247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_779_im = _RAND_1248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_780_re = _RAND_1249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_780_im = _RAND_1250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_781_re = _RAND_1251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  _T_781_im = _RAND_1252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  _T_782_re = _RAND_1253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  _T_782_im = _RAND_1254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  _T_783_re = _RAND_1255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  _T_783_im = _RAND_1256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  _T_784_re = _RAND_1257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  _T_784_im = _RAND_1258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  _T_785_re = _RAND_1259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  _T_785_im = _RAND_1260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  _T_786_re = _RAND_1261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  _T_786_im = _RAND_1262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  _T_787_re = _RAND_1263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  _T_787_im = _RAND_1264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  _T_788_re = _RAND_1265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  _T_788_im = _RAND_1266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  _T_789_re = _RAND_1267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  _T_789_im = _RAND_1268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  _T_790_re = _RAND_1269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  _T_790_im = _RAND_1270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  _T_791_re = _RAND_1271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  _T_791_im = _RAND_1272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  _T_792_re = _RAND_1273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  _T_792_im = _RAND_1274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  _T_793_re = _RAND_1275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  _T_793_im = _RAND_1276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  _T_794_re = _RAND_1277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  _T_794_im = _RAND_1278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  _T_795_re = _RAND_1279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  _T_795_im = _RAND_1280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  _T_797_re = _RAND_1281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  _T_797_im = _RAND_1282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  _T_798_re = _RAND_1283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  _T_798_im = _RAND_1284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  _T_799_re = _RAND_1285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  _T_799_im = _RAND_1286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  _T_800_re = _RAND_1287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  _T_800_im = _RAND_1288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  _T_801_re = _RAND_1289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  _T_801_im = _RAND_1290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  _T_802_re = _RAND_1291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  _T_802_im = _RAND_1292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  _T_803_re = _RAND_1293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  _T_803_im = _RAND_1294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  _T_804_re = _RAND_1295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  _T_804_im = _RAND_1296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  _T_805_re = _RAND_1297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  _T_805_im = _RAND_1298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  _T_806_re = _RAND_1299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  _T_806_im = _RAND_1300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  _T_807_re = _RAND_1301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  _T_807_im = _RAND_1302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  _T_808_re = _RAND_1303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  _T_808_im = _RAND_1304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  _T_809_re = _RAND_1305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  _T_809_im = _RAND_1306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  _T_810_re = _RAND_1307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  _T_810_im = _RAND_1308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  _T_811_re = _RAND_1309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  _T_811_im = _RAND_1310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  _T_812_re = _RAND_1311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  _T_812_im = _RAND_1312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  _T_813_re = _RAND_1313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  _T_813_im = _RAND_1314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  _T_814_re = _RAND_1315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  _T_814_im = _RAND_1316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  _T_815_re = _RAND_1317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  _T_815_im = _RAND_1318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  _T_816_re = _RAND_1319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  _T_816_im = _RAND_1320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  _T_817_re = _RAND_1321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  _T_817_im = _RAND_1322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  _T_818_re = _RAND_1323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  _T_818_im = _RAND_1324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  _T_819_re = _RAND_1325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  _T_819_im = _RAND_1326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  _T_820_re = _RAND_1327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  _T_820_im = _RAND_1328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  _T_821_re = _RAND_1329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  _T_821_im = _RAND_1330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  _T_822_re = _RAND_1331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  _T_822_im = _RAND_1332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  _T_823_re = _RAND_1333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  _T_823_im = _RAND_1334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  _T_824_re = _RAND_1335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  _T_824_im = _RAND_1336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  _T_825_re = _RAND_1337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  _T_825_im = _RAND_1338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  _T_826_re = _RAND_1339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  _T_826_im = _RAND_1340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  _T_827_re = _RAND_1341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  _T_827_im = _RAND_1342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  _T_828_re = _RAND_1343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  _T_828_im = _RAND_1344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  _T_833_re = _RAND_1345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  _T_833_im = _RAND_1346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  _T_834_re = _RAND_1347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  _T_834_im = _RAND_1348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  _T_835_re = _RAND_1349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  _T_835_im = _RAND_1350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  _T_836_re = _RAND_1351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  _T_836_im = _RAND_1352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  _T_837_re = _RAND_1353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  _T_837_im = _RAND_1354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  _T_838_re = _RAND_1355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  _T_838_im = _RAND_1356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  _T_839_re = _RAND_1357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  _T_839_im = _RAND_1358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  _T_840_re = _RAND_1359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  _T_840_im = _RAND_1360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  _T_841_re = _RAND_1361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  _T_841_im = _RAND_1362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  _T_842_re = _RAND_1363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  _T_842_im = _RAND_1364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  _T_843_re = _RAND_1365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  _T_843_im = _RAND_1366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  _T_844_re = _RAND_1367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  _T_844_im = _RAND_1368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  _T_845_re = _RAND_1369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  _T_845_im = _RAND_1370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  _T_846_re = _RAND_1371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  _T_846_im = _RAND_1372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  _T_847_re = _RAND_1373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  _T_847_im = _RAND_1374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  _T_848_re = _RAND_1375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  _T_848_im = _RAND_1376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  _T_849_re = _RAND_1377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  _T_849_im = _RAND_1378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  _T_850_re = _RAND_1379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  _T_850_im = _RAND_1380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  _T_851_re = _RAND_1381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  _T_851_im = _RAND_1382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  _T_852_re = _RAND_1383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  _T_852_im = _RAND_1384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  _T_853_re = _RAND_1385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  _T_853_im = _RAND_1386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  _T_854_re = _RAND_1387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  _T_854_im = _RAND_1388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  _T_855_re = _RAND_1389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  _T_855_im = _RAND_1390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  _T_856_re = _RAND_1391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  _T_856_im = _RAND_1392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  _T_857_re = _RAND_1393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  _T_857_im = _RAND_1394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  _T_858_re = _RAND_1395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  _T_858_im = _RAND_1396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  _T_859_re = _RAND_1397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  _T_859_im = _RAND_1398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  _T_860_re = _RAND_1399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  _T_860_im = _RAND_1400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  _T_861_re = _RAND_1401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  _T_861_im = _RAND_1402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  _T_862_re = _RAND_1403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  _T_862_im = _RAND_1404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  _T_863_re = _RAND_1405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  _T_863_im = _RAND_1406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  _T_864_re = _RAND_1407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  _T_864_im = _RAND_1408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  _T_866_re = _RAND_1409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  _T_866_im = _RAND_1410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  _T_867_re = _RAND_1411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  _T_867_im = _RAND_1412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  _T_868_re = _RAND_1413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  _T_868_im = _RAND_1414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  _T_869_re = _RAND_1415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  _T_869_im = _RAND_1416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  _T_870_re = _RAND_1417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  _T_870_im = _RAND_1418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  _T_871_re = _RAND_1419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  _T_871_im = _RAND_1420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  _T_872_re = _RAND_1421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  _T_872_im = _RAND_1422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  _T_873_re = _RAND_1423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  _T_873_im = _RAND_1424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  _T_874_re = _RAND_1425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  _T_874_im = _RAND_1426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  _T_875_re = _RAND_1427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  _T_875_im = _RAND_1428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  _T_876_re = _RAND_1429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  _T_876_im = _RAND_1430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  _T_877_re = _RAND_1431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  _T_877_im = _RAND_1432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  _T_878_re = _RAND_1433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  _T_878_im = _RAND_1434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  _T_879_re = _RAND_1435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  _T_879_im = _RAND_1436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  _T_880_re = _RAND_1437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  _T_880_im = _RAND_1438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  _T_881_re = _RAND_1439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  _T_881_im = _RAND_1440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  _T_886_re = _RAND_1441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  _T_886_im = _RAND_1442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  _T_887_re = _RAND_1443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  _T_887_im = _RAND_1444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  _T_888_re = _RAND_1445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  _T_888_im = _RAND_1446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  _T_889_re = _RAND_1447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  _T_889_im = _RAND_1448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  _T_890_re = _RAND_1449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  _T_890_im = _RAND_1450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  _T_891_re = _RAND_1451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  _T_891_im = _RAND_1452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  _T_892_re = _RAND_1453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  _T_892_im = _RAND_1454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  _T_893_re = _RAND_1455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  _T_893_im = _RAND_1456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  _T_894_re = _RAND_1457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  _T_894_im = _RAND_1458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  _T_895_re = _RAND_1459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  _T_895_im = _RAND_1460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  _T_896_re = _RAND_1461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  _T_896_im = _RAND_1462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  _T_897_re = _RAND_1463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  _T_897_im = _RAND_1464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  _T_898_re = _RAND_1465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  _T_898_im = _RAND_1466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  _T_899_re = _RAND_1467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  _T_899_im = _RAND_1468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  _T_900_re = _RAND_1469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  _T_900_im = _RAND_1470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  _T_901_re = _RAND_1471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  _T_901_im = _RAND_1472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  _T_903_re = _RAND_1473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  _T_903_im = _RAND_1474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  _T_904_re = _RAND_1475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  _T_904_im = _RAND_1476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  _T_905_re = _RAND_1477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  _T_905_im = _RAND_1478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  _T_906_re = _RAND_1479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  _T_906_im = _RAND_1480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  _T_907_re = _RAND_1481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  _T_907_im = _RAND_1482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  _T_908_re = _RAND_1483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  _T_908_im = _RAND_1484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  _T_909_re = _RAND_1485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  _T_909_im = _RAND_1486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  _T_910_re = _RAND_1487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  _T_910_im = _RAND_1488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  _T_915_re = _RAND_1489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  _T_915_im = _RAND_1490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  _T_916_re = _RAND_1491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  _T_916_im = _RAND_1492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  _T_917_re = _RAND_1493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  _T_917_im = _RAND_1494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  _T_918_re = _RAND_1495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  _T_918_im = _RAND_1496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  _T_919_re = _RAND_1497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  _T_919_im = _RAND_1498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  _T_920_re = _RAND_1499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  _T_920_im = _RAND_1500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  _T_921_re = _RAND_1501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  _T_921_im = _RAND_1502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  _T_922_re = _RAND_1503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  _T_922_im = _RAND_1504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  _T_924_re = _RAND_1505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  _T_924_im = _RAND_1506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  _T_925_re = _RAND_1507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  _T_925_im = _RAND_1508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  _T_926_re = _RAND_1509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  _T_926_im = _RAND_1510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  _T_927_re = _RAND_1511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  _T_927_im = _RAND_1512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  _T_932_re = _RAND_1513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  _T_932_im = _RAND_1514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  _T_933_re = _RAND_1515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  _T_933_im = _RAND_1516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  _T_934_re = _RAND_1517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  _T_934_im = _RAND_1518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  _T_935_re = _RAND_1519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  _T_935_im = _RAND_1520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  _T_937_re = _RAND_1521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  _T_937_im = _RAND_1522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  _T_938_re = _RAND_1523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  _T_938_im = _RAND_1524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  _T_943_re = _RAND_1525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  _T_943_im = _RAND_1526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  _T_944_re = _RAND_1527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  _T_944_im = _RAND_1528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  _T_946_re = _RAND_1529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  _T_946_im = _RAND_1530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  out1D1_re = _RAND_1531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  out1D1_im = _RAND_1532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  _T_947_re = _RAND_1533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  _T_947_im = _RAND_1534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  _T_948_re = _RAND_1535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  _T_948_im = _RAND_1536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  _T_949 = _RAND_1537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  _T_950 = _RAND_1538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  _T_951 = _RAND_1539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  _T_952 = _RAND_1540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  _T_953 = _RAND_1541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  _T_954 = _RAND_1542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1543 = {1{`RANDOM}};
  _T_955 = _RAND_1543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1544 = {1{`RANDOM}};
  _T_956 = _RAND_1544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1545 = {1{`RANDOM}};
  _T_957 = _RAND_1545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1546 = {1{`RANDOM}};
  _T_958 = _RAND_1546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1547 = {1{`RANDOM}};
  _T_959 = _RAND_1547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1548 = {1{`RANDOM}};
  _T_960 = _RAND_1548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1549 = {1{`RANDOM}};
  _T_961 = _RAND_1549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1550 = {1{`RANDOM}};
  _T_962 = _RAND_1550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1551 = {1{`RANDOM}};
  _T_963 = _RAND_1551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1552 = {1{`RANDOM}};
  _T_964 = _RAND_1552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1553 = {1{`RANDOM}};
  _T_965 = _RAND_1553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1554 = {1{`RANDOM}};
  _T_966 = _RAND_1554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1555 = {1{`RANDOM}};
  _T_967 = _RAND_1555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1556 = {1{`RANDOM}};
  _T_968 = _RAND_1556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1557 = {1{`RANDOM}};
  _T_969 = _RAND_1557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1558 = {1{`RANDOM}};
  _T_970 = _RAND_1558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1559 = {1{`RANDOM}};
  _T_971 = _RAND_1559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1560 = {1{`RANDOM}};
  _T_972 = _RAND_1560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1561 = {1{`RANDOM}};
  _T_973 = _RAND_1561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1562 = {1{`RANDOM}};
  _T_974 = _RAND_1562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1563 = {1{`RANDOM}};
  _T_975 = _RAND_1563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1564 = {1{`RANDOM}};
  _T_976 = _RAND_1564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1565 = {1{`RANDOM}};
  _T_977 = _RAND_1565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1566 = {1{`RANDOM}};
  _T_978 = _RAND_1566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1567 = {1{`RANDOM}};
  _T_979 = _RAND_1567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1568 = {1{`RANDOM}};
  _T_980 = _RAND_1568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1569 = {1{`RANDOM}};
  _T_981 = _RAND_1569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1570 = {1{`RANDOM}};
  _T_982 = _RAND_1570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1571 = {1{`RANDOM}};
  _T_983 = _RAND_1571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1572 = {1{`RANDOM}};
  _T_984 = _RAND_1572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1573 = {1{`RANDOM}};
  _T_985 = _RAND_1573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1574 = {1{`RANDOM}};
  _T_986 = _RAND_1574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1575 = {1{`RANDOM}};
  _T_987 = _RAND_1575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1576 = {1{`RANDOM}};
  _T_988 = _RAND_1576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1577 = {1{`RANDOM}};
  _T_989 = _RAND_1577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1578 = {1{`RANDOM}};
  _T_990 = _RAND_1578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1579 = {1{`RANDOM}};
  _T_991 = _RAND_1579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1580 = {1{`RANDOM}};
  _T_992 = _RAND_1580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1581 = {1{`RANDOM}};
  _T_993 = _RAND_1581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1582 = {1{`RANDOM}};
  _T_994 = _RAND_1582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1583 = {1{`RANDOM}};
  _T_995 = _RAND_1583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1584 = {1{`RANDOM}};
  _T_996 = _RAND_1584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1585 = {1{`RANDOM}};
  _T_997 = _RAND_1585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1586 = {1{`RANDOM}};
  _T_998 = _RAND_1586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1587 = {1{`RANDOM}};
  _T_999 = _RAND_1587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1588 = {1{`RANDOM}};
  _T_1000 = _RAND_1588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1589 = {1{`RANDOM}};
  _T_1001 = _RAND_1589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1590 = {1{`RANDOM}};
  _T_1002 = _RAND_1590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1591 = {1{`RANDOM}};
  _T_1003 = _RAND_1591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1592 = {1{`RANDOM}};
  _T_1004 = _RAND_1592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1593 = {1{`RANDOM}};
  _T_1005 = _RAND_1593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1594 = {1{`RANDOM}};
  _T_1006 = _RAND_1594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1595 = {1{`RANDOM}};
  _T_1007 = _RAND_1595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1596 = {1{`RANDOM}};
  _T_1008 = _RAND_1596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1597 = {1{`RANDOM}};
  _T_1009 = _RAND_1597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1598 = {1{`RANDOM}};
  _T_1010 = _RAND_1598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1599 = {1{`RANDOM}};
  _T_1011 = _RAND_1599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1600 = {1{`RANDOM}};
  _T_1012 = _RAND_1600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1601 = {1{`RANDOM}};
  _T_1013 = _RAND_1601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1602 = {1{`RANDOM}};
  _T_1014 = _RAND_1602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1603 = {1{`RANDOM}};
  _T_1015 = _RAND_1603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1604 = {1{`RANDOM}};
  _T_1016 = _RAND_1604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1605 = {1{`RANDOM}};
  _T_1017 = _RAND_1605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1606 = {1{`RANDOM}};
  _T_1018 = _RAND_1606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1607 = {1{`RANDOM}};
  _T_1019 = _RAND_1607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1608 = {1{`RANDOM}};
  _T_1020 = _RAND_1608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1609 = {1{`RANDOM}};
  _T_1021 = _RAND_1609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1610 = {1{`RANDOM}};
  _T_1022 = _RAND_1610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1611 = {1{`RANDOM}};
  _T_1023 = _RAND_1611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1612 = {1{`RANDOM}};
  _T_1024 = _RAND_1612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1613 = {1{`RANDOM}};
  _T_1025 = _RAND_1613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1614 = {1{`RANDOM}};
  _T_1026 = _RAND_1614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1615 = {1{`RANDOM}};
  _T_1027 = _RAND_1615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1616 = {1{`RANDOM}};
  _T_1028 = _RAND_1616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1617 = {1{`RANDOM}};
  _T_1029 = _RAND_1617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1618 = {1{`RANDOM}};
  _T_1030 = _RAND_1618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1619 = {1{`RANDOM}};
  _T_1031 = _RAND_1619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1620 = {1{`RANDOM}};
  _T_1032 = _RAND_1620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1621 = {1{`RANDOM}};
  _T_1033 = _RAND_1621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1622 = {1{`RANDOM}};
  _T_1034 = _RAND_1622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1623 = {1{`RANDOM}};
  _T_1035 = _RAND_1623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1624 = {1{`RANDOM}};
  _T_1036 = _RAND_1624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1625 = {1{`RANDOM}};
  _T_1037 = _RAND_1625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1626 = {1{`RANDOM}};
  _T_1038 = _RAND_1626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1627 = {1{`RANDOM}};
  _T_1039 = _RAND_1627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1628 = {1{`RANDOM}};
  _T_1040 = _RAND_1628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1629 = {1{`RANDOM}};
  _T_1041 = _RAND_1629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1630 = {1{`RANDOM}};
  _T_1042 = _RAND_1630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1631 = {1{`RANDOM}};
  _T_1043 = _RAND_1631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1632 = {1{`RANDOM}};
  _T_1044 = _RAND_1632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1633 = {1{`RANDOM}};
  _T_1045 = _RAND_1633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1634 = {1{`RANDOM}};
  _T_1046 = _RAND_1634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1635 = {1{`RANDOM}};
  _T_1047 = _RAND_1635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1636 = {1{`RANDOM}};
  _T_1048 = _RAND_1636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1637 = {1{`RANDOM}};
  _T_1049 = _RAND_1637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1638 = {1{`RANDOM}};
  _T_1050 = _RAND_1638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1639 = {1{`RANDOM}};
  _T_1051 = _RAND_1639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1640 = {1{`RANDOM}};
  _T_1052 = _RAND_1640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1641 = {1{`RANDOM}};
  _T_1053 = _RAND_1641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1642 = {1{`RANDOM}};
  _T_1054 = _RAND_1642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1643 = {1{`RANDOM}};
  _T_1055 = _RAND_1643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1644 = {1{`RANDOM}};
  _T_1056 = _RAND_1644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1645 = {1{`RANDOM}};
  _T_1057 = _RAND_1645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1646 = {1{`RANDOM}};
  _T_1058 = _RAND_1646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1647 = {1{`RANDOM}};
  _T_1059 = _RAND_1647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1648 = {1{`RANDOM}};
  _T_1060 = _RAND_1648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1649 = {1{`RANDOM}};
  _T_1061 = _RAND_1649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1650 = {1{`RANDOM}};
  _T_1062 = _RAND_1650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1651 = {1{`RANDOM}};
  _T_1063 = _RAND_1651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1652 = {1{`RANDOM}};
  _T_1064 = _RAND_1652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1653 = {1{`RANDOM}};
  _T_1065 = _RAND_1653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1654 = {1{`RANDOM}};
  _T_1066 = _RAND_1654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1655 = {1{`RANDOM}};
  _T_1067 = _RAND_1655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1656 = {1{`RANDOM}};
  _T_1068 = _RAND_1656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1657 = {1{`RANDOM}};
  _T_1069 = _RAND_1657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1658 = {1{`RANDOM}};
  _T_1070 = _RAND_1658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1659 = {1{`RANDOM}};
  _T_1071 = _RAND_1659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1660 = {1{`RANDOM}};
  _T_1072 = _RAND_1660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1661 = {1{`RANDOM}};
  _T_1073 = _RAND_1661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1662 = {1{`RANDOM}};
  _T_1074 = _RAND_1662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1663 = {1{`RANDOM}};
  _T_1075 = _RAND_1663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1664 = {1{`RANDOM}};
  _T_1076 = _RAND_1664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1665 = {1{`RANDOM}};
  _T_1077 = _RAND_1665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1666 = {1{`RANDOM}};
  _T_1078 = _RAND_1666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1667 = {1{`RANDOM}};
  _T_1079 = _RAND_1667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1668 = {1{`RANDOM}};
  _T_1080 = _RAND_1668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1669 = {1{`RANDOM}};
  _T_1081 = _RAND_1669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1670 = {1{`RANDOM}};
  _T_1082 = _RAND_1670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1671 = {1{`RANDOM}};
  _T_1083 = _RAND_1671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1672 = {1{`RANDOM}};
  _T_1084 = _RAND_1672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1673 = {1{`RANDOM}};
  _T_1085 = _RAND_1673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1674 = {1{`RANDOM}};
  _T_1086 = _RAND_1674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1675 = {1{`RANDOM}};
  _T_1087 = _RAND_1675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1676 = {1{`RANDOM}};
  _T_1088 = _RAND_1676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1677 = {1{`RANDOM}};
  _T_1089 = _RAND_1677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1678 = {1{`RANDOM}};
  _T_1090 = _RAND_1678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1679 = {1{`RANDOM}};
  _T_1091 = _RAND_1679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1680 = {1{`RANDOM}};
  _T_1092 = _RAND_1680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1681 = {1{`RANDOM}};
  _T_1093 = _RAND_1681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1682 = {1{`RANDOM}};
  _T_1094 = _RAND_1682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1683 = {1{`RANDOM}};
  _T_1095 = _RAND_1683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1684 = {1{`RANDOM}};
  _T_1096 = _RAND_1684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1685 = {1{`RANDOM}};
  _T_1097 = _RAND_1685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1686 = {1{`RANDOM}};
  _T_1098 = _RAND_1686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1687 = {1{`RANDOM}};
  _T_1099 = _RAND_1687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1688 = {1{`RANDOM}};
  _T_1100 = _RAND_1688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1689 = {1{`RANDOM}};
  _T_1101 = _RAND_1689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1690 = {1{`RANDOM}};
  _T_1102 = _RAND_1690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1691 = {1{`RANDOM}};
  _T_1103 = _RAND_1691[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1692 = {1{`RANDOM}};
  _T_1104 = _RAND_1692[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1693 = {1{`RANDOM}};
  _T_1105 = _RAND_1693[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1694 = {1{`RANDOM}};
  _T_1106 = _RAND_1694[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1695 = {1{`RANDOM}};
  _T_1107 = _RAND_1695[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1696 = {1{`RANDOM}};
  _T_1108 = _RAND_1696[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1697 = {1{`RANDOM}};
  _T_1109 = _RAND_1697[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1698 = {1{`RANDOM}};
  _T_1110 = _RAND_1698[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1699 = {1{`RANDOM}};
  _T_1111 = _RAND_1699[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1700 = {1{`RANDOM}};
  _T_1112 = _RAND_1700[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1701 = {1{`RANDOM}};
  _T_1113 = _RAND_1701[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1702 = {1{`RANDOM}};
  _T_1114 = _RAND_1702[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1703 = {1{`RANDOM}};
  _T_1115 = _RAND_1703[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1704 = {1{`RANDOM}};
  _T_1116 = _RAND_1704[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1705 = {1{`RANDOM}};
  _T_1117 = _RAND_1705[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1706 = {1{`RANDOM}};
  _T_1118 = _RAND_1706[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1707 = {1{`RANDOM}};
  _T_1119 = _RAND_1707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1708 = {1{`RANDOM}};
  _T_1120 = _RAND_1708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1709 = {1{`RANDOM}};
  _T_1121 = _RAND_1709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1710 = {1{`RANDOM}};
  _T_1122 = _RAND_1710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1711 = {1{`RANDOM}};
  _T_1123 = _RAND_1711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1712 = {1{`RANDOM}};
  _T_1124 = _RAND_1712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1713 = {1{`RANDOM}};
  _T_1125 = _RAND_1713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1714 = {1{`RANDOM}};
  _T_1126 = _RAND_1714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1715 = {1{`RANDOM}};
  _T_1127 = _RAND_1715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1716 = {1{`RANDOM}};
  _T_1128 = _RAND_1716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1717 = {1{`RANDOM}};
  _T_1129 = _RAND_1717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1718 = {1{`RANDOM}};
  _T_1130 = _RAND_1718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1719 = {1{`RANDOM}};
  _T_1131 = _RAND_1719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1720 = {1{`RANDOM}};
  _T_1132 = _RAND_1720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1721 = {1{`RANDOM}};
  _T_1133 = _RAND_1721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1722 = {1{`RANDOM}};
  _T_1134 = _RAND_1722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1723 = {1{`RANDOM}};
  _T_1135 = _RAND_1723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1724 = {1{`RANDOM}};
  _T_1136 = _RAND_1724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1725 = {1{`RANDOM}};
  _T_1137 = _RAND_1725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1726 = {1{`RANDOM}};
  _T_1138 = _RAND_1726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1727 = {1{`RANDOM}};
  _T_1139 = _RAND_1727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1728 = {1{`RANDOM}};
  _T_1140 = _RAND_1728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1729 = {1{`RANDOM}};
  _T_1141 = _RAND_1729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1730 = {1{`RANDOM}};
  _T_1142 = _RAND_1730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1731 = {1{`RANDOM}};
  _T_1143 = _RAND_1731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1732 = {1{`RANDOM}};
  _T_1144 = _RAND_1732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1733 = {1{`RANDOM}};
  _T_1145 = _RAND_1733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1734 = {1{`RANDOM}};
  _T_1146 = _RAND_1734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1735 = {1{`RANDOM}};
  _T_1147 = _RAND_1735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1736 = {1{`RANDOM}};
  _T_1148 = _RAND_1736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1737 = {1{`RANDOM}};
  _T_1149 = _RAND_1737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1738 = {1{`RANDOM}};
  _T_1150 = _RAND_1738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1739 = {1{`RANDOM}};
  _T_1151 = _RAND_1739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1740 = {1{`RANDOM}};
  _T_1152 = _RAND_1740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1741 = {1{`RANDOM}};
  _T_1153 = _RAND_1741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1742 = {1{`RANDOM}};
  _T_1154 = _RAND_1742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1743 = {1{`RANDOM}};
  _T_1155 = _RAND_1743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1744 = {1{`RANDOM}};
  _T_1156 = _RAND_1744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1745 = {1{`RANDOM}};
  _T_1157 = _RAND_1745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1746 = {1{`RANDOM}};
  _T_1158 = _RAND_1746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1747 = {1{`RANDOM}};
  _T_1159 = _RAND_1747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1748 = {1{`RANDOM}};
  _T_1160 = _RAND_1748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1749 = {1{`RANDOM}};
  _T_1161 = _RAND_1749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1750 = {1{`RANDOM}};
  _T_1162 = _RAND_1750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1751 = {1{`RANDOM}};
  _T_1163 = _RAND_1751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1752 = {1{`RANDOM}};
  _T_1164 = _RAND_1752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1753 = {1{`RANDOM}};
  _T_1165 = _RAND_1753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1754 = {1{`RANDOM}};
  _T_1166 = _RAND_1754[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1755 = {1{`RANDOM}};
  _T_1167 = _RAND_1755[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1756 = {1{`RANDOM}};
  _T_1168 = _RAND_1756[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1757 = {1{`RANDOM}};
  _T_1169 = _RAND_1757[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1758 = {1{`RANDOM}};
  _T_1170 = _RAND_1758[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1759 = {1{`RANDOM}};
  _T_1171 = _RAND_1759[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1760 = {1{`RANDOM}};
  _T_1172 = _RAND_1760[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1761 = {1{`RANDOM}};
  _T_1173 = _RAND_1761[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1762 = {1{`RANDOM}};
  _T_1174 = _RAND_1762[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1763 = {1{`RANDOM}};
  _T_1175 = _RAND_1763[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1764 = {1{`RANDOM}};
  _T_1176 = _RAND_1764[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1765 = {1{`RANDOM}};
  _T_1177 = _RAND_1765[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1766 = {1{`RANDOM}};
  _T_1178 = _RAND_1766[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1767 = {1{`RANDOM}};
  _T_1179 = _RAND_1767[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1768 = {1{`RANDOM}};
  _T_1180 = _RAND_1768[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1769 = {1{`RANDOM}};
  _T_1181 = _RAND_1769[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1770 = {1{`RANDOM}};
  _T_1182 = _RAND_1770[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1771 = {1{`RANDOM}};
  _T_1183 = _RAND_1771[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1772 = {1{`RANDOM}};
  _T_1184 = _RAND_1772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1773 = {1{`RANDOM}};
  _T_1185 = _RAND_1773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1774 = {1{`RANDOM}};
  _T_1186 = _RAND_1774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1775 = {1{`RANDOM}};
  _T_1187 = _RAND_1775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1776 = {1{`RANDOM}};
  _T_1188 = _RAND_1776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1777 = {1{`RANDOM}};
  _T_1189 = _RAND_1777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1778 = {1{`RANDOM}};
  _T_1190 = _RAND_1778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1779 = {1{`RANDOM}};
  _T_1191 = _RAND_1779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1780 = {1{`RANDOM}};
  _T_1192 = _RAND_1780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1781 = {1{`RANDOM}};
  _T_1193 = _RAND_1781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1782 = {1{`RANDOM}};
  _T_1194 = _RAND_1782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1783 = {1{`RANDOM}};
  _T_1195 = _RAND_1783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1784 = {1{`RANDOM}};
  _T_1196 = _RAND_1784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1785 = {1{`RANDOM}};
  _T_1197 = _RAND_1785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1786 = {1{`RANDOM}};
  _T_1198 = _RAND_1786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1787 = {1{`RANDOM}};
  _T_1199 = _RAND_1787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1788 = {1{`RANDOM}};
  _T_1200 = _RAND_1788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1789 = {1{`RANDOM}};
  _T_1201 = _RAND_1789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1790 = {1{`RANDOM}};
  _T_1202 = _RAND_1790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1791 = {1{`RANDOM}};
  _T_1203 = _RAND_1791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1792 = {1{`RANDOM}};
  _T_1204 = _RAND_1792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1793 = {1{`RANDOM}};
  _T_1205 = _RAND_1793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1794 = {1{`RANDOM}};
  _T_1206 = _RAND_1794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1795 = {1{`RANDOM}};
  _T_1207 = _RAND_1795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1796 = {1{`RANDOM}};
  _T_1208 = _RAND_1796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1797 = {1{`RANDOM}};
  _T_1209 = _RAND_1797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1798 = {1{`RANDOM}};
  _T_1210 = _RAND_1798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1799 = {1{`RANDOM}};
  _T_1211 = _RAND_1799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1800 = {1{`RANDOM}};
  _T_1212 = _RAND_1800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1801 = {1{`RANDOM}};
  _T_1213 = _RAND_1801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1802 = {1{`RANDOM}};
  _T_1214 = _RAND_1802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1803 = {1{`RANDOM}};
  _T_1215 = _RAND_1803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1804 = {1{`RANDOM}};
  _T_1216 = _RAND_1804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1805 = {1{`RANDOM}};
  _T_1217 = _RAND_1805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1806 = {1{`RANDOM}};
  _T_1218 = _RAND_1806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1807 = {1{`RANDOM}};
  _T_1219 = _RAND_1807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1808 = {1{`RANDOM}};
  _T_1220 = _RAND_1808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1809 = {1{`RANDOM}};
  _T_1221 = _RAND_1809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1810 = {1{`RANDOM}};
  _T_1222 = _RAND_1810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1811 = {1{`RANDOM}};
  _T_1223 = _RAND_1811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1812 = {1{`RANDOM}};
  _T_1224 = _RAND_1812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1813 = {1{`RANDOM}};
  _T_1225 = _RAND_1813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1814 = {1{`RANDOM}};
  _T_1226 = _RAND_1814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1815 = {1{`RANDOM}};
  _T_1227 = _RAND_1815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1816 = {1{`RANDOM}};
  _T_1228 = _RAND_1816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1817 = {1{`RANDOM}};
  _T_1229 = _RAND_1817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1818 = {1{`RANDOM}};
  _T_1230 = _RAND_1818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1819 = {1{`RANDOM}};
  _T_1231 = _RAND_1819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1820 = {1{`RANDOM}};
  _T_1232 = _RAND_1820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1821 = {1{`RANDOM}};
  _T_1233 = _RAND_1821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1822 = {1{`RANDOM}};
  _T_1234 = _RAND_1822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1823 = {1{`RANDOM}};
  _T_1235 = _RAND_1823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1824 = {1{`RANDOM}};
  _T_1236 = _RAND_1824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1825 = {1{`RANDOM}};
  _T_1237 = _RAND_1825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1826 = {1{`RANDOM}};
  _T_1238 = _RAND_1826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1827 = {1{`RANDOM}};
  _T_1239 = _RAND_1827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1828 = {1{`RANDOM}};
  _T_1240 = _RAND_1828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1829 = {1{`RANDOM}};
  _T_1241 = _RAND_1829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1830 = {1{`RANDOM}};
  _T_1242 = _RAND_1830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1831 = {1{`RANDOM}};
  _T_1243 = _RAND_1831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1832 = {1{`RANDOM}};
  _T_1244 = _RAND_1832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1833 = {1{`RANDOM}};
  _T_1245 = _RAND_1833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1834 = {1{`RANDOM}};
  _T_1246 = _RAND_1834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1835 = {1{`RANDOM}};
  _T_1247 = _RAND_1835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1836 = {1{`RANDOM}};
  _T_1248 = _RAND_1836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1837 = {1{`RANDOM}};
  _T_1249 = _RAND_1837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1838 = {1{`RANDOM}};
  _T_1250 = _RAND_1838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1839 = {1{`RANDOM}};
  _T_1251 = _RAND_1839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1840 = {1{`RANDOM}};
  _T_1252 = _RAND_1840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1841 = {1{`RANDOM}};
  _T_1253 = _RAND_1841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1842 = {1{`RANDOM}};
  _T_1254 = _RAND_1842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1843 = {1{`RANDOM}};
  _T_1255 = _RAND_1843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1844 = {1{`RANDOM}};
  _T_1256 = _RAND_1844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1845 = {1{`RANDOM}};
  _T_1257 = _RAND_1845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1846 = {1{`RANDOM}};
  _T_1258 = _RAND_1846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1847 = {1{`RANDOM}};
  _T_1259 = _RAND_1847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1848 = {1{`RANDOM}};
  _T_1260 = _RAND_1848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1849 = {1{`RANDOM}};
  _T_1261 = _RAND_1849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1850 = {1{`RANDOM}};
  _T_1262 = _RAND_1850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1851 = {1{`RANDOM}};
  _T_1263 = _RAND_1851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1852 = {1{`RANDOM}};
  _T_1264 = _RAND_1852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1853 = {1{`RANDOM}};
  _T_1265 = _RAND_1853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1854 = {1{`RANDOM}};
  _T_1266 = _RAND_1854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1855 = {1{`RANDOM}};
  _T_1267 = _RAND_1855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1856 = {1{`RANDOM}};
  _T_1268 = _RAND_1856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1857 = {1{`RANDOM}};
  _T_1269 = _RAND_1857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1858 = {1{`RANDOM}};
  _T_1270 = _RAND_1858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1859 = {1{`RANDOM}};
  _T_1271 = _RAND_1859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1860 = {1{`RANDOM}};
  _T_1272 = _RAND_1860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1861 = {1{`RANDOM}};
  _T_1273 = _RAND_1861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1862 = {1{`RANDOM}};
  _T_1274 = _RAND_1862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1863 = {1{`RANDOM}};
  _T_1275 = _RAND_1863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1864 = {1{`RANDOM}};
  _T_1276 = _RAND_1864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1865 = {1{`RANDOM}};
  _T_1277 = _RAND_1865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1866 = {1{`RANDOM}};
  _T_1278 = _RAND_1866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1867 = {1{`RANDOM}};
  _T_1279 = _RAND_1867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1868 = {1{`RANDOM}};
  _T_1280 = _RAND_1868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1869 = {1{`RANDOM}};
  _T_1281 = _RAND_1869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1870 = {1{`RANDOM}};
  _T_1282 = _RAND_1870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1871 = {1{`RANDOM}};
  _T_1283 = _RAND_1871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1872 = {1{`RANDOM}};
  _T_1284 = _RAND_1872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1873 = {1{`RANDOM}};
  _T_1285 = _RAND_1873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1874 = {1{`RANDOM}};
  _T_1286 = _RAND_1874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1875 = {1{`RANDOM}};
  _T_1287 = _RAND_1875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1876 = {1{`RANDOM}};
  _T_1288 = _RAND_1876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1877 = {1{`RANDOM}};
  _T_1289 = _RAND_1877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1878 = {1{`RANDOM}};
  _T_1290 = _RAND_1878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1879 = {1{`RANDOM}};
  _T_1291 = _RAND_1879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1880 = {1{`RANDOM}};
  _T_1292 = _RAND_1880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1881 = {1{`RANDOM}};
  _T_1293 = _RAND_1881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1882 = {1{`RANDOM}};
  _T_1294 = _RAND_1882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1883 = {1{`RANDOM}};
  _T_1295 = _RAND_1883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1884 = {1{`RANDOM}};
  _T_1296 = _RAND_1884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1885 = {1{`RANDOM}};
  _T_1297 = _RAND_1885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1886 = {1{`RANDOM}};
  _T_1298 = _RAND_1886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1887 = {1{`RANDOM}};
  _T_1299 = _RAND_1887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1888 = {1{`RANDOM}};
  _T_1300 = _RAND_1888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1889 = {1{`RANDOM}};
  _T_1301 = _RAND_1889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1890 = {1{`RANDOM}};
  _T_1302 = _RAND_1890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1891 = {1{`RANDOM}};
  _T_1303 = _RAND_1891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1892 = {1{`RANDOM}};
  _T_1304 = _RAND_1892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1893 = {1{`RANDOM}};
  _T_1305 = _RAND_1893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1894 = {1{`RANDOM}};
  _T_1306 = _RAND_1894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1895 = {1{`RANDOM}};
  _T_1307 = _RAND_1895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1896 = {1{`RANDOM}};
  _T_1308 = _RAND_1896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1897 = {1{`RANDOM}};
  _T_1309 = _RAND_1897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1898 = {1{`RANDOM}};
  _T_1310 = _RAND_1898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1899 = {1{`RANDOM}};
  _T_1311 = _RAND_1899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1900 = {1{`RANDOM}};
  _T_1312 = _RAND_1900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1901 = {1{`RANDOM}};
  _T_1313 = _RAND_1901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1902 = {1{`RANDOM}};
  _T_1314 = _RAND_1902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1903 = {1{`RANDOM}};
  _T_1315 = _RAND_1903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1904 = {1{`RANDOM}};
  _T_1316 = _RAND_1904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1905 = {1{`RANDOM}};
  _T_1317 = _RAND_1905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1906 = {1{`RANDOM}};
  _T_1318 = _RAND_1906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1907 = {1{`RANDOM}};
  _T_1319 = _RAND_1907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1908 = {1{`RANDOM}};
  _T_1320 = _RAND_1908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1909 = {1{`RANDOM}};
  _T_1321 = _RAND_1909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1910 = {1{`RANDOM}};
  _T_1322 = _RAND_1910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1911 = {1{`RANDOM}};
  _T_1323 = _RAND_1911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1912 = {1{`RANDOM}};
  _T_1324 = _RAND_1912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1913 = {1{`RANDOM}};
  _T_1325 = _RAND_1913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1914 = {1{`RANDOM}};
  _T_1326 = _RAND_1914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1915 = {1{`RANDOM}};
  _T_1327 = _RAND_1915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1916 = {1{`RANDOM}};
  _T_1328 = _RAND_1916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1917 = {1{`RANDOM}};
  _T_1329 = _RAND_1917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1918 = {1{`RANDOM}};
  _T_1330 = _RAND_1918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1919 = {1{`RANDOM}};
  _T_1331 = _RAND_1919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1920 = {1{`RANDOM}};
  _T_1332 = _RAND_1920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1921 = {1{`RANDOM}};
  _T_1333 = _RAND_1921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1922 = {1{`RANDOM}};
  _T_1334 = _RAND_1922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1923 = {1{`RANDOM}};
  _T_1335 = _RAND_1923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1924 = {1{`RANDOM}};
  _T_1336 = _RAND_1924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1925 = {1{`RANDOM}};
  _T_1337 = _RAND_1925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1926 = {1{`RANDOM}};
  _T_1338 = _RAND_1926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1927 = {1{`RANDOM}};
  _T_1339 = _RAND_1927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1928 = {1{`RANDOM}};
  _T_1340 = _RAND_1928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1929 = {1{`RANDOM}};
  _T_1341 = _RAND_1929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1930 = {1{`RANDOM}};
  _T_1342 = _RAND_1930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1931 = {1{`RANDOM}};
  _T_1343 = _RAND_1931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1932 = {1{`RANDOM}};
  _T_1344 = _RAND_1932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1933 = {1{`RANDOM}};
  _T_1345 = _RAND_1933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1934 = {1{`RANDOM}};
  _T_1346 = _RAND_1934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1935 = {1{`RANDOM}};
  _T_1347 = _RAND_1935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1936 = {1{`RANDOM}};
  _T_1348 = _RAND_1936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1937 = {1{`RANDOM}};
  _T_1349 = _RAND_1937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1938 = {1{`RANDOM}};
  _T_1350 = _RAND_1938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1939 = {1{`RANDOM}};
  _T_1351 = _RAND_1939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1940 = {1{`RANDOM}};
  _T_1352 = _RAND_1940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1941 = {1{`RANDOM}};
  _T_1353 = _RAND_1941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1942 = {1{`RANDOM}};
  _T_1354 = _RAND_1942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1943 = {1{`RANDOM}};
  _T_1355 = _RAND_1943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1944 = {1{`RANDOM}};
  _T_1356 = _RAND_1944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1945 = {1{`RANDOM}};
  _T_1357 = _RAND_1945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1946 = {1{`RANDOM}};
  _T_1358 = _RAND_1946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1947 = {1{`RANDOM}};
  _T_1359 = _RAND_1947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1948 = {1{`RANDOM}};
  _T_1360 = _RAND_1948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1949 = {1{`RANDOM}};
  _T_1361 = _RAND_1949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1950 = {1{`RANDOM}};
  _T_1362 = _RAND_1950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1951 = {1{`RANDOM}};
  _T_1363 = _RAND_1951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1952 = {1{`RANDOM}};
  _T_1364 = _RAND_1952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1953 = {1{`RANDOM}};
  _T_1365 = _RAND_1953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1954 = {1{`RANDOM}};
  _T_1366 = _RAND_1954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1955 = {1{`RANDOM}};
  _T_1367 = _RAND_1955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1956 = {1{`RANDOM}};
  _T_1368 = _RAND_1956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1957 = {1{`RANDOM}};
  _T_1369 = _RAND_1957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1958 = {1{`RANDOM}};
  _T_1370 = _RAND_1958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1959 = {1{`RANDOM}};
  _T_1371 = _RAND_1959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1960 = {1{`RANDOM}};
  _T_1372 = _RAND_1960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1961 = {1{`RANDOM}};
  _T_1373 = _RAND_1961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1962 = {1{`RANDOM}};
  _T_1374 = _RAND_1962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1963 = {1{`RANDOM}};
  _T_1375 = _RAND_1963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1964 = {1{`RANDOM}};
  _T_1376 = _RAND_1964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1965 = {1{`RANDOM}};
  _T_1377 = _RAND_1965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1966 = {1{`RANDOM}};
  _T_1378 = _RAND_1966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1967 = {1{`RANDOM}};
  _T_1379 = _RAND_1967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1968 = {1{`RANDOM}};
  _T_1380 = _RAND_1968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1969 = {1{`RANDOM}};
  _T_1381 = _RAND_1969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1970 = {1{`RANDOM}};
  _T_1382 = _RAND_1970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1971 = {1{`RANDOM}};
  _T_1383 = _RAND_1971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1972 = {1{`RANDOM}};
  _T_1384 = _RAND_1972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1973 = {1{`RANDOM}};
  _T_1385 = _RAND_1973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1974 = {1{`RANDOM}};
  _T_1386 = _RAND_1974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1975 = {1{`RANDOM}};
  _T_1387 = _RAND_1975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1976 = {1{`RANDOM}};
  _T_1388 = _RAND_1976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1977 = {1{`RANDOM}};
  _T_1389 = _RAND_1977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1978 = {1{`RANDOM}};
  _T_1390 = _RAND_1978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1979 = {1{`RANDOM}};
  _T_1391 = _RAND_1979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1980 = {1{`RANDOM}};
  _T_1392 = _RAND_1980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1981 = {1{`RANDOM}};
  _T_1393 = _RAND_1981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1982 = {1{`RANDOM}};
  _T_1394 = _RAND_1982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1983 = {1{`RANDOM}};
  _T_1395 = _RAND_1983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1984 = {1{`RANDOM}};
  _T_1396 = _RAND_1984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1985 = {1{`RANDOM}};
  _T_1397 = _RAND_1985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1986 = {1{`RANDOM}};
  _T_1398 = _RAND_1986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1987 = {1{`RANDOM}};
  _T_1399 = _RAND_1987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1988 = {1{`RANDOM}};
  _T_1400 = _RAND_1988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1989 = {1{`RANDOM}};
  _T_1401 = _RAND_1989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1990 = {1{`RANDOM}};
  _T_1402 = _RAND_1990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1991 = {1{`RANDOM}};
  _T_1403 = _RAND_1991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1992 = {1{`RANDOM}};
  _T_1404 = _RAND_1992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1993 = {1{`RANDOM}};
  _T_1405 = _RAND_1993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1994 = {1{`RANDOM}};
  _T_1406 = _RAND_1994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1995 = {1{`RANDOM}};
  _T_1407 = _RAND_1995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1996 = {1{`RANDOM}};
  _T_1408 = _RAND_1996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1997 = {1{`RANDOM}};
  _T_1409 = _RAND_1997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1998 = {1{`RANDOM}};
  _T_1410 = _RAND_1998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1999 = {1{`RANDOM}};
  _T_1411 = _RAND_1999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2000 = {1{`RANDOM}};
  _T_1412 = _RAND_2000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2001 = {1{`RANDOM}};
  _T_1413 = _RAND_2001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2002 = {1{`RANDOM}};
  _T_1414 = _RAND_2002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2003 = {1{`RANDOM}};
  _T_1415 = _RAND_2003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2004 = {1{`RANDOM}};
  _T_1416 = _RAND_2004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2005 = {1{`RANDOM}};
  _T_1417 = _RAND_2005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2006 = {1{`RANDOM}};
  _T_1418 = _RAND_2006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2007 = {1{`RANDOM}};
  _T_1419 = _RAND_2007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2008 = {1{`RANDOM}};
  _T_1420 = _RAND_2008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2009 = {1{`RANDOM}};
  _T_1421 = _RAND_2009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2010 = {1{`RANDOM}};
  _T_1422 = _RAND_2010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2011 = {1{`RANDOM}};
  _T_1423 = _RAND_2011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2012 = {1{`RANDOM}};
  _T_1424 = _RAND_2012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2013 = {1{`RANDOM}};
  _T_1425 = _RAND_2013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2014 = {1{`RANDOM}};
  _T_1426 = _RAND_2014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2015 = {1{`RANDOM}};
  _T_1427 = _RAND_2015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2016 = {1{`RANDOM}};
  _T_1428 = _RAND_2016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2017 = {1{`RANDOM}};
  _T_1429 = _RAND_2017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2018 = {1{`RANDOM}};
  _T_1430 = _RAND_2018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2019 = {1{`RANDOM}};
  _T_1431 = _RAND_2019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2020 = {1{`RANDOM}};
  _T_1432 = _RAND_2020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2021 = {1{`RANDOM}};
  _T_1433 = _RAND_2021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2022 = {1{`RANDOM}};
  _T_1434 = _RAND_2022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2023 = {1{`RANDOM}};
  _T_1435 = _RAND_2023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2024 = {1{`RANDOM}};
  _T_1436 = _RAND_2024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2025 = {1{`RANDOM}};
  _T_1437 = _RAND_2025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2026 = {1{`RANDOM}};
  _T_1438 = _RAND_2026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2027 = {1{`RANDOM}};
  _T_1439 = _RAND_2027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2028 = {1{`RANDOM}};
  _T_1440 = _RAND_2028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2029 = {1{`RANDOM}};
  _T_1441 = _RAND_2029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2030 = {1{`RANDOM}};
  _T_1442 = _RAND_2030[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2031 = {1{`RANDOM}};
  _T_1443 = _RAND_2031[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2032 = {1{`RANDOM}};
  _T_1444 = _RAND_2032[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2033 = {1{`RANDOM}};
  _T_1445 = _RAND_2033[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2034 = {1{`RANDOM}};
  _T_1446 = _RAND_2034[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2035 = {1{`RANDOM}};
  _T_1447 = _RAND_2035[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2036 = {1{`RANDOM}};
  _T_1448 = _RAND_2036[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2037 = {1{`RANDOM}};
  _T_1449 = _RAND_2037[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2038 = {1{`RANDOM}};
  _T_1450 = _RAND_2038[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2039 = {1{`RANDOM}};
  _T_1451 = _RAND_2039[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2040 = {1{`RANDOM}};
  _T_1452 = _RAND_2040[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2041 = {1{`RANDOM}};
  _T_1453 = _RAND_2041[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2042 = {1{`RANDOM}};
  _T_1454 = _RAND_2042[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2043 = {1{`RANDOM}};
  _T_1455 = _RAND_2043[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2044 = {1{`RANDOM}};
  _T_1456 = _RAND_2044[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2045 = {1{`RANDOM}};
  _T_1457 = _RAND_2045[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2046 = {1{`RANDOM}};
  _T_1458 = _RAND_2046[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2047 = {1{`RANDOM}};
  _T_1459 = _RAND_2047[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2048 = {1{`RANDOM}};
  _T_1460 = _RAND_2048[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 9'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    _T_146_re <= io_dIn_re;
    _T_146_im <= io_dIn_im;
    _T_147_re <= _T_146_re;
    _T_147_im <= _T_146_im;
    _T_148_re <= _T_147_re;
    _T_148_im <= _T_147_im;
    _T_149_re <= _T_148_re;
    _T_149_im <= _T_148_im;
    _T_150_re <= _T_149_re;
    _T_150_im <= _T_149_im;
    _T_151_re <= _T_150_re;
    _T_151_im <= _T_150_im;
    _T_152_re <= _T_151_re;
    _T_152_im <= _T_151_im;
    _T_153_re <= _T_152_re;
    _T_153_im <= _T_152_im;
    _T_154_re <= _T_153_re;
    _T_154_im <= _T_153_im;
    _T_155_re <= _T_154_re;
    _T_155_im <= _T_154_im;
    _T_156_re <= _T_155_re;
    _T_156_im <= _T_155_im;
    _T_157_re <= _T_156_re;
    _T_157_im <= _T_156_im;
    _T_158_re <= _T_157_re;
    _T_158_im <= _T_157_im;
    _T_159_re <= _T_158_re;
    _T_159_im <= _T_158_im;
    _T_160_re <= _T_159_re;
    _T_160_im <= _T_159_im;
    _T_161_re <= _T_160_re;
    _T_161_im <= _T_160_im;
    _T_162_re <= _T_161_re;
    _T_162_im <= _T_161_im;
    _T_163_re <= _T_162_re;
    _T_163_im <= _T_162_im;
    _T_164_re <= _T_163_re;
    _T_164_im <= _T_163_im;
    _T_165_re <= _T_164_re;
    _T_165_im <= _T_164_im;
    _T_166_re <= _T_165_re;
    _T_166_im <= _T_165_im;
    _T_167_re <= _T_166_re;
    _T_167_im <= _T_166_im;
    _T_168_re <= _T_167_re;
    _T_168_im <= _T_167_im;
    _T_169_re <= _T_168_re;
    _T_169_im <= _T_168_im;
    _T_170_re <= _T_169_re;
    _T_170_im <= _T_169_im;
    _T_171_re <= _T_170_re;
    _T_171_im <= _T_170_im;
    _T_172_re <= _T_171_re;
    _T_172_im <= _T_171_im;
    _T_173_re <= _T_172_re;
    _T_173_im <= _T_172_im;
    _T_174_re <= _T_173_re;
    _T_174_im <= _T_173_im;
    _T_175_re <= _T_174_re;
    _T_175_im <= _T_174_im;
    _T_176_re <= _T_175_re;
    _T_176_im <= _T_175_im;
    _T_177_re <= _T_176_re;
    _T_177_im <= _T_176_im;
    _T_178_re <= _T_177_re;
    _T_178_im <= _T_177_im;
    _T_179_re <= _T_178_re;
    _T_179_im <= _T_178_im;
    _T_180_re <= _T_179_re;
    _T_180_im <= _T_179_im;
    _T_181_re <= _T_180_re;
    _T_181_im <= _T_180_im;
    _T_182_re <= _T_181_re;
    _T_182_im <= _T_181_im;
    _T_183_re <= _T_182_re;
    _T_183_im <= _T_182_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_325_re <= _T_324_re;
    _T_325_im <= _T_324_im;
    _T_326_re <= _T_325_re;
    _T_326_im <= _T_325_im;
    _T_327_re <= _T_326_re;
    _T_327_im <= _T_326_im;
    _T_328_re <= _T_327_re;
    _T_328_im <= _T_327_im;
    _T_329_re <= _T_328_re;
    _T_329_im <= _T_328_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_393_re <= _T_392_re;
    _T_393_im <= _T_392_im;
    _T_394_re <= _T_393_re;
    _T_394_im <= _T_393_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_403_re <= Butterfly_io_out2_re;
    _T_403_im <= Butterfly_io_out2_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_406_re <= _T_405_re;
    _T_406_im <= _T_405_im;
    _T_407_re <= _T_406_re;
    _T_407_im <= _T_406_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_409_re <= _T_408_re;
    _T_409_im <= _T_408_im;
    _T_410_re <= _T_409_re;
    _T_410_im <= _T_409_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_535_re <= Switch_io_out1_re;
    _T_535_im <= Switch_io_out1_im;
    _T_536_re <= _T_535_re;
    _T_536_im <= _T_535_im;
    _T_537_re <= _T_536_re;
    _T_537_im <= _T_536_im;
    _T_538_re <= _T_537_re;
    _T_538_im <= _T_537_im;
    _T_539_re <= _T_538_re;
    _T_539_im <= _T_538_im;
    _T_540_re <= _T_539_re;
    _T_540_im <= _T_539_im;
    _T_541_re <= _T_540_re;
    _T_541_im <= _T_540_im;
    _T_542_re <= _T_541_re;
    _T_542_im <= _T_541_im;
    _T_543_re <= _T_542_re;
    _T_543_im <= _T_542_im;
    _T_544_re <= _T_543_re;
    _T_544_im <= _T_543_im;
    _T_545_re <= _T_544_re;
    _T_545_im <= _T_544_im;
    _T_546_re <= _T_545_re;
    _T_546_im <= _T_545_im;
    _T_547_re <= _T_546_re;
    _T_547_im <= _T_546_im;
    _T_548_re <= _T_547_re;
    _T_548_im <= _T_547_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_664_re <= Butterfly_1_io_out2_re;
    _T_664_im <= Butterfly_1_io_out2_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_671_re <= _T_670_re;
    _T_671_im <= _T_670_im;
    _T_672_re <= _T_671_re;
    _T_672_im <= _T_671_im;
    _T_673_re <= _T_672_re;
    _T_673_im <= _T_672_im;
    _T_674_re <= _T_673_re;
    _T_674_im <= _T_673_im;
    _T_675_re <= _T_674_re;
    _T_675_im <= _T_674_im;
    _T_676_re <= _T_675_re;
    _T_676_im <= _T_675_im;
    _T_677_re <= _T_676_re;
    _T_677_im <= _T_676_im;
    _T_678_re <= _T_677_re;
    _T_678_im <= _T_677_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_732_re <= Switch_1_io_out1_re;
    _T_732_im <= Switch_1_io_out1_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_736_re <= _T_735_re;
    _T_736_im <= _T_735_im;
    _T_737_re <= _T_736_re;
    _T_737_im <= _T_736_im;
    _T_738_re <= _T_737_re;
    _T_738_im <= _T_737_im;
    _T_739_re <= _T_738_re;
    _T_739_im <= _T_738_im;
    _T_740_re <= _T_739_re;
    _T_740_im <= _T_739_im;
    _T_741_re <= _T_740_re;
    _T_741_im <= _T_740_im;
    _T_742_re <= _T_741_re;
    _T_742_im <= _T_741_im;
    _T_743_re <= _T_742_re;
    _T_743_im <= _T_742_im;
    _T_744_re <= _T_743_re;
    _T_744_im <= _T_743_im;
    _T_745_re <= _T_744_re;
    _T_745_im <= _T_744_im;
    _T_746_re <= _T_745_re;
    _T_746_im <= _T_745_im;
    _T_747_re <= _T_746_re;
    _T_747_im <= _T_746_im;
    _T_748_re <= _T_747_re;
    _T_748_im <= _T_747_im;
    _T_749_re <= _T_748_re;
    _T_749_im <= _T_748_im;
    _T_750_re <= _T_749_re;
    _T_750_im <= _T_749_im;
    _T_751_re <= _T_750_re;
    _T_751_im <= _T_750_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_797_re <= Butterfly_2_io_out2_re;
    _T_797_im <= Butterfly_2_io_out2_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_808_re <= _T_807_re;
    _T_808_im <= _T_807_im;
    _T_809_re <= _T_808_re;
    _T_809_im <= _T_808_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_811_re <= _T_810_re;
    _T_811_im <= _T_810_im;
    _T_812_re <= _T_811_re;
    _T_812_im <= _T_811_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_815_re <= _T_814_re;
    _T_815_im <= _T_814_im;
    _T_816_re <= _T_815_re;
    _T_816_im <= _T_815_im;
    _T_817_re <= _T_816_re;
    _T_817_im <= _T_816_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_833_re <= Switch_2_io_out1_re;
    _T_833_im <= Switch_2_io_out1_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_841_re <= _T_840_re;
    _T_841_im <= _T_840_im;
    _T_842_re <= _T_841_re;
    _T_842_im <= _T_841_im;
    _T_843_re <= _T_842_re;
    _T_843_im <= _T_842_im;
    _T_844_re <= _T_843_re;
    _T_844_im <= _T_843_im;
    _T_845_re <= _T_844_re;
    _T_845_im <= _T_844_im;
    _T_846_re <= _T_845_re;
    _T_846_im <= _T_845_im;
    _T_847_re <= _T_846_re;
    _T_847_im <= _T_846_im;
    _T_848_re <= _T_847_re;
    _T_848_im <= _T_847_im;
    _T_849_re <= _T_848_re;
    _T_849_im <= _T_848_im;
    _T_850_re <= _T_849_re;
    _T_850_im <= _T_849_im;
    _T_851_re <= _T_850_re;
    _T_851_im <= _T_850_im;
    _T_852_re <= _T_851_re;
    _T_852_im <= _T_851_im;
    _T_853_re <= _T_852_re;
    _T_853_im <= _T_852_im;
    _T_854_re <= _T_853_re;
    _T_854_im <= _T_853_im;
    _T_855_re <= _T_854_re;
    _T_855_im <= _T_854_im;
    _T_856_re <= _T_855_re;
    _T_856_im <= _T_855_im;
    _T_857_re <= _T_856_re;
    _T_857_im <= _T_856_im;
    _T_858_re <= _T_857_re;
    _T_858_im <= _T_857_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_866_re <= Butterfly_3_io_out2_re;
    _T_866_im <= Butterfly_3_io_out2_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_881_re <= _T_880_re;
    _T_881_im <= _T_880_im;
    _T_886_re <= Switch_3_io_out1_re;
    _T_886_im <= Switch_3_io_out1_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_890_re <= _T_889_re;
    _T_890_im <= _T_889_im;
    _T_891_re <= _T_890_re;
    _T_891_im <= _T_890_im;
    _T_892_re <= _T_891_re;
    _T_892_im <= _T_891_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_898_re <= _T_897_re;
    _T_898_im <= _T_897_im;
    _T_899_re <= _T_898_re;
    _T_899_im <= _T_898_im;
    _T_900_re <= _T_899_re;
    _T_900_im <= _T_899_im;
    _T_901_re <= _T_900_re;
    _T_901_im <= _T_900_im;
    _T_903_re <= Butterfly_4_io_out2_re;
    _T_903_im <= Butterfly_4_io_out2_im;
    _T_904_re <= _T_903_re;
    _T_904_im <= _T_903_im;
    _T_905_re <= _T_904_re;
    _T_905_im <= _T_904_im;
    _T_906_re <= _T_905_re;
    _T_906_im <= _T_905_im;
    _T_907_re <= _T_906_re;
    _T_907_im <= _T_906_im;
    _T_908_re <= _T_907_re;
    _T_908_im <= _T_907_im;
    _T_909_re <= _T_908_re;
    _T_909_im <= _T_908_im;
    _T_910_re <= _T_909_re;
    _T_910_im <= _T_909_im;
    _T_915_re <= Switch_4_io_out1_re;
    _T_915_im <= Switch_4_io_out1_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_922_re <= _T_921_re;
    _T_922_im <= _T_921_im;
    _T_924_re <= Butterfly_5_io_out2_re;
    _T_924_im <= Butterfly_5_io_out2_im;
    _T_925_re <= _T_924_re;
    _T_925_im <= _T_924_im;
    _T_926_re <= _T_925_re;
    _T_926_im <= _T_925_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_932_re <= Switch_5_io_out1_re;
    _T_932_im <= Switch_5_io_out1_im;
    _T_933_re <= _T_932_re;
    _T_933_im <= _T_932_im;
    _T_934_re <= _T_933_re;
    _T_934_im <= _T_933_im;
    _T_935_re <= _T_934_re;
    _T_935_im <= _T_934_im;
    _T_937_re <= Butterfly_6_io_out2_re;
    _T_937_im <= Butterfly_6_io_out2_im;
    _T_938_re <= _T_937_re;
    _T_938_im <= _T_937_im;
    _T_943_re <= Switch_6_io_out1_re;
    _T_943_im <= Switch_6_io_out1_im;
    _T_944_re <= _T_943_re;
    _T_944_im <= _T_943_im;
    _T_946_re <= Butterfly_7_io_out2_re;
    _T_946_im <= Butterfly_7_io_out2_im;
    out1D1_re <= Switch_7_io_out1_re;
    out1D1_im <= Switch_7_io_out1_im;
    _T_947_re <= ComplexAdd_io_res_re;
    _T_947_im <= ComplexAdd_io_res_im;
    _T_948_re <= ComplexSub_io_res_re;
    _T_948_im <= ComplexSub_io_res_im;
    _T_949 <= io_din_valid;
    _T_950 <= _T_949;
    _T_951 <= _T_950;
    _T_952 <= _T_951;
    _T_953 <= _T_952;
    _T_954 <= _T_953;
    _T_955 <= _T_954;
    _T_956 <= _T_955;
    _T_957 <= _T_956;
    _T_958 <= _T_957;
    _T_959 <= _T_958;
    _T_960 <= _T_959;
    _T_961 <= _T_960;
    _T_962 <= _T_961;
    _T_963 <= _T_962;
    _T_964 <= _T_963;
    _T_965 <= _T_964;
    _T_966 <= _T_965;
    _T_967 <= _T_966;
    _T_968 <= _T_967;
    _T_969 <= _T_968;
    _T_970 <= _T_969;
    _T_971 <= _T_970;
    _T_972 <= _T_971;
    _T_973 <= _T_972;
    _T_974 <= _T_973;
    _T_975 <= _T_974;
    _T_976 <= _T_975;
    _T_977 <= _T_976;
    _T_978 <= _T_977;
    _T_979 <= _T_978;
    _T_980 <= _T_979;
    _T_981 <= _T_980;
    _T_982 <= _T_981;
    _T_983 <= _T_982;
    _T_984 <= _T_983;
    _T_985 <= _T_984;
    _T_986 <= _T_985;
    _T_987 <= _T_986;
    _T_988 <= _T_987;
    _T_989 <= _T_988;
    _T_990 <= _T_989;
    _T_991 <= _T_990;
    _T_992 <= _T_991;
    _T_993 <= _T_992;
    _T_994 <= _T_993;
    _T_995 <= _T_994;
    _T_996 <= _T_995;
    _T_997 <= _T_996;
    _T_998 <= _T_997;
    _T_999 <= _T_998;
    _T_1000 <= _T_999;
    _T_1001 <= _T_1000;
    _T_1002 <= _T_1001;
    _T_1003 <= _T_1002;
    _T_1004 <= _T_1003;
    _T_1005 <= _T_1004;
    _T_1006 <= _T_1005;
    _T_1007 <= _T_1006;
    _T_1008 <= _T_1007;
    _T_1009 <= _T_1008;
    _T_1010 <= _T_1009;
    _T_1011 <= _T_1010;
    _T_1012 <= _T_1011;
    _T_1013 <= _T_1012;
    _T_1014 <= _T_1013;
    _T_1015 <= _T_1014;
    _T_1016 <= _T_1015;
    _T_1017 <= _T_1016;
    _T_1018 <= _T_1017;
    _T_1019 <= _T_1018;
    _T_1020 <= _T_1019;
    _T_1021 <= _T_1020;
    _T_1022 <= _T_1021;
    _T_1023 <= _T_1022;
    _T_1024 <= _T_1023;
    _T_1025 <= _T_1024;
    _T_1026 <= _T_1025;
    _T_1027 <= _T_1026;
    _T_1028 <= _T_1027;
    _T_1029 <= _T_1028;
    _T_1030 <= _T_1029;
    _T_1031 <= _T_1030;
    _T_1032 <= _T_1031;
    _T_1033 <= _T_1032;
    _T_1034 <= _T_1033;
    _T_1035 <= _T_1034;
    _T_1036 <= _T_1035;
    _T_1037 <= _T_1036;
    _T_1038 <= _T_1037;
    _T_1039 <= _T_1038;
    _T_1040 <= _T_1039;
    _T_1041 <= _T_1040;
    _T_1042 <= _T_1041;
    _T_1043 <= _T_1042;
    _T_1044 <= _T_1043;
    _T_1045 <= _T_1044;
    _T_1046 <= _T_1045;
    _T_1047 <= _T_1046;
    _T_1048 <= _T_1047;
    _T_1049 <= _T_1048;
    _T_1050 <= _T_1049;
    _T_1051 <= _T_1050;
    _T_1052 <= _T_1051;
    _T_1053 <= _T_1052;
    _T_1054 <= _T_1053;
    _T_1055 <= _T_1054;
    _T_1056 <= _T_1055;
    _T_1057 <= _T_1056;
    _T_1058 <= _T_1057;
    _T_1059 <= _T_1058;
    _T_1060 <= _T_1059;
    _T_1061 <= _T_1060;
    _T_1062 <= _T_1061;
    _T_1063 <= _T_1062;
    _T_1064 <= _T_1063;
    _T_1065 <= _T_1064;
    _T_1066 <= _T_1065;
    _T_1067 <= _T_1066;
    _T_1068 <= _T_1067;
    _T_1069 <= _T_1068;
    _T_1070 <= _T_1069;
    _T_1071 <= _T_1070;
    _T_1072 <= _T_1071;
    _T_1073 <= _T_1072;
    _T_1074 <= _T_1073;
    _T_1075 <= _T_1074;
    _T_1076 <= _T_1075;
    _T_1077 <= _T_1076;
    _T_1078 <= _T_1077;
    _T_1079 <= _T_1078;
    _T_1080 <= _T_1079;
    _T_1081 <= _T_1080;
    _T_1082 <= _T_1081;
    _T_1083 <= _T_1082;
    _T_1084 <= _T_1083;
    _T_1085 <= _T_1084;
    _T_1086 <= _T_1085;
    _T_1087 <= _T_1086;
    _T_1088 <= _T_1087;
    _T_1089 <= _T_1088;
    _T_1090 <= _T_1089;
    _T_1091 <= _T_1090;
    _T_1092 <= _T_1091;
    _T_1093 <= _T_1092;
    _T_1094 <= _T_1093;
    _T_1095 <= _T_1094;
    _T_1096 <= _T_1095;
    _T_1097 <= _T_1096;
    _T_1098 <= _T_1097;
    _T_1099 <= _T_1098;
    _T_1100 <= _T_1099;
    _T_1101 <= _T_1100;
    _T_1102 <= _T_1101;
    _T_1103 <= _T_1102;
    _T_1104 <= _T_1103;
    _T_1105 <= _T_1104;
    _T_1106 <= _T_1105;
    _T_1107 <= _T_1106;
    _T_1108 <= _T_1107;
    _T_1109 <= _T_1108;
    _T_1110 <= _T_1109;
    _T_1111 <= _T_1110;
    _T_1112 <= _T_1111;
    _T_1113 <= _T_1112;
    _T_1114 <= _T_1113;
    _T_1115 <= _T_1114;
    _T_1116 <= _T_1115;
    _T_1117 <= _T_1116;
    _T_1118 <= _T_1117;
    _T_1119 <= _T_1118;
    _T_1120 <= _T_1119;
    _T_1121 <= _T_1120;
    _T_1122 <= _T_1121;
    _T_1123 <= _T_1122;
    _T_1124 <= _T_1123;
    _T_1125 <= _T_1124;
    _T_1126 <= _T_1125;
    _T_1127 <= _T_1126;
    _T_1128 <= _T_1127;
    _T_1129 <= _T_1128;
    _T_1130 <= _T_1129;
    _T_1131 <= _T_1130;
    _T_1132 <= _T_1131;
    _T_1133 <= _T_1132;
    _T_1134 <= _T_1133;
    _T_1135 <= _T_1134;
    _T_1136 <= _T_1135;
    _T_1137 <= _T_1136;
    _T_1138 <= _T_1137;
    _T_1139 <= _T_1138;
    _T_1140 <= _T_1139;
    _T_1141 <= _T_1140;
    _T_1142 <= _T_1141;
    _T_1143 <= _T_1142;
    _T_1144 <= _T_1143;
    _T_1145 <= _T_1144;
    _T_1146 <= _T_1145;
    _T_1147 <= _T_1146;
    _T_1148 <= _T_1147;
    _T_1149 <= _T_1148;
    _T_1150 <= _T_1149;
    _T_1151 <= _T_1150;
    _T_1152 <= _T_1151;
    _T_1153 <= _T_1152;
    _T_1154 <= _T_1153;
    _T_1155 <= _T_1154;
    _T_1156 <= _T_1155;
    _T_1157 <= _T_1156;
    _T_1158 <= _T_1157;
    _T_1159 <= _T_1158;
    _T_1160 <= _T_1159;
    _T_1161 <= _T_1160;
    _T_1162 <= _T_1161;
    _T_1163 <= _T_1162;
    _T_1164 <= _T_1163;
    _T_1165 <= _T_1164;
    _T_1166 <= _T_1165;
    _T_1167 <= _T_1166;
    _T_1168 <= _T_1167;
    _T_1169 <= _T_1168;
    _T_1170 <= _T_1169;
    _T_1171 <= _T_1170;
    _T_1172 <= _T_1171;
    _T_1173 <= _T_1172;
    _T_1174 <= _T_1173;
    _T_1175 <= _T_1174;
    _T_1176 <= _T_1175;
    _T_1177 <= _T_1176;
    _T_1178 <= _T_1177;
    _T_1179 <= _T_1178;
    _T_1180 <= _T_1179;
    _T_1181 <= _T_1180;
    _T_1182 <= _T_1181;
    _T_1183 <= _T_1182;
    _T_1184 <= _T_1183;
    _T_1185 <= _T_1184;
    _T_1186 <= _T_1185;
    _T_1187 <= _T_1186;
    _T_1188 <= _T_1187;
    _T_1189 <= _T_1188;
    _T_1190 <= _T_1189;
    _T_1191 <= _T_1190;
    _T_1192 <= _T_1191;
    _T_1193 <= _T_1192;
    _T_1194 <= _T_1193;
    _T_1195 <= _T_1194;
    _T_1196 <= _T_1195;
    _T_1197 <= _T_1196;
    _T_1198 <= _T_1197;
    _T_1199 <= _T_1198;
    _T_1200 <= _T_1199;
    _T_1201 <= _T_1200;
    _T_1202 <= _T_1201;
    _T_1203 <= _T_1202;
    _T_1204 <= _T_1203;
    _T_1205 <= _T_1204;
    _T_1206 <= _T_1205;
    _T_1207 <= _T_1206;
    _T_1208 <= _T_1207;
    _T_1209 <= _T_1208;
    _T_1210 <= _T_1209;
    _T_1211 <= _T_1210;
    _T_1212 <= _T_1211;
    _T_1213 <= _T_1212;
    _T_1214 <= _T_1213;
    _T_1215 <= _T_1214;
    _T_1216 <= _T_1215;
    _T_1217 <= _T_1216;
    _T_1218 <= _T_1217;
    _T_1219 <= _T_1218;
    _T_1220 <= _T_1219;
    _T_1221 <= _T_1220;
    _T_1222 <= _T_1221;
    _T_1223 <= _T_1222;
    _T_1224 <= _T_1223;
    _T_1225 <= _T_1224;
    _T_1226 <= _T_1225;
    _T_1227 <= _T_1226;
    _T_1228 <= _T_1227;
    _T_1229 <= _T_1228;
    _T_1230 <= _T_1229;
    _T_1231 <= _T_1230;
    _T_1232 <= _T_1231;
    _T_1233 <= _T_1232;
    _T_1234 <= _T_1233;
    _T_1235 <= _T_1234;
    _T_1236 <= _T_1235;
    _T_1237 <= _T_1236;
    _T_1238 <= _T_1237;
    _T_1239 <= _T_1238;
    _T_1240 <= _T_1239;
    _T_1241 <= _T_1240;
    _T_1242 <= _T_1241;
    _T_1243 <= _T_1242;
    _T_1244 <= _T_1243;
    _T_1245 <= _T_1244;
    _T_1246 <= _T_1245;
    _T_1247 <= _T_1246;
    _T_1248 <= _T_1247;
    _T_1249 <= _T_1248;
    _T_1250 <= _T_1249;
    _T_1251 <= _T_1250;
    _T_1252 <= _T_1251;
    _T_1253 <= _T_1252;
    _T_1254 <= _T_1253;
    _T_1255 <= _T_1254;
    _T_1256 <= _T_1255;
    _T_1257 <= _T_1256;
    _T_1258 <= _T_1257;
    _T_1259 <= _T_1258;
    _T_1260 <= _T_1259;
    _T_1261 <= _T_1260;
    _T_1262 <= _T_1261;
    _T_1263 <= _T_1262;
    _T_1264 <= _T_1263;
    _T_1265 <= _T_1264;
    _T_1266 <= _T_1265;
    _T_1267 <= _T_1266;
    _T_1268 <= _T_1267;
    _T_1269 <= _T_1268;
    _T_1270 <= _T_1269;
    _T_1271 <= _T_1270;
    _T_1272 <= _T_1271;
    _T_1273 <= _T_1272;
    _T_1274 <= _T_1273;
    _T_1275 <= _T_1274;
    _T_1276 <= _T_1275;
    _T_1277 <= _T_1276;
    _T_1278 <= _T_1277;
    _T_1279 <= _T_1278;
    _T_1280 <= _T_1279;
    _T_1281 <= _T_1280;
    _T_1282 <= _T_1281;
    _T_1283 <= _T_1282;
    _T_1284 <= _T_1283;
    _T_1285 <= _T_1284;
    _T_1286 <= _T_1285;
    _T_1287 <= _T_1286;
    _T_1288 <= _T_1287;
    _T_1289 <= _T_1288;
    _T_1290 <= _T_1289;
    _T_1291 <= _T_1290;
    _T_1292 <= _T_1291;
    _T_1293 <= _T_1292;
    _T_1294 <= _T_1293;
    _T_1295 <= _T_1294;
    _T_1296 <= _T_1295;
    _T_1297 <= _T_1296;
    _T_1298 <= _T_1297;
    _T_1299 <= _T_1298;
    _T_1300 <= _T_1299;
    _T_1301 <= _T_1300;
    _T_1302 <= _T_1301;
    _T_1303 <= _T_1302;
    _T_1304 <= _T_1303;
    _T_1305 <= _T_1304;
    _T_1306 <= _T_1305;
    _T_1307 <= _T_1306;
    _T_1308 <= _T_1307;
    _T_1309 <= _T_1308;
    _T_1310 <= _T_1309;
    _T_1311 <= _T_1310;
    _T_1312 <= _T_1311;
    _T_1313 <= _T_1312;
    _T_1314 <= _T_1313;
    _T_1315 <= _T_1314;
    _T_1316 <= _T_1315;
    _T_1317 <= _T_1316;
    _T_1318 <= _T_1317;
    _T_1319 <= _T_1318;
    _T_1320 <= _T_1319;
    _T_1321 <= _T_1320;
    _T_1322 <= _T_1321;
    _T_1323 <= _T_1322;
    _T_1324 <= _T_1323;
    _T_1325 <= _T_1324;
    _T_1326 <= _T_1325;
    _T_1327 <= _T_1326;
    _T_1328 <= _T_1327;
    _T_1329 <= _T_1328;
    _T_1330 <= _T_1329;
    _T_1331 <= _T_1330;
    _T_1332 <= _T_1331;
    _T_1333 <= _T_1332;
    _T_1334 <= _T_1333;
    _T_1335 <= _T_1334;
    _T_1336 <= _T_1335;
    _T_1337 <= _T_1336;
    _T_1338 <= _T_1337;
    _T_1339 <= _T_1338;
    _T_1340 <= _T_1339;
    _T_1341 <= _T_1340;
    _T_1342 <= _T_1341;
    _T_1343 <= _T_1342;
    _T_1344 <= _T_1343;
    _T_1345 <= _T_1344;
    _T_1346 <= _T_1345;
    _T_1347 <= _T_1346;
    _T_1348 <= _T_1347;
    _T_1349 <= _T_1348;
    _T_1350 <= _T_1349;
    _T_1351 <= _T_1350;
    _T_1352 <= _T_1351;
    _T_1353 <= _T_1352;
    _T_1354 <= _T_1353;
    _T_1355 <= _T_1354;
    _T_1356 <= _T_1355;
    _T_1357 <= _T_1356;
    _T_1358 <= _T_1357;
    _T_1359 <= _T_1358;
    _T_1360 <= _T_1359;
    _T_1361 <= _T_1360;
    _T_1362 <= _T_1361;
    _T_1363 <= _T_1362;
    _T_1364 <= _T_1363;
    _T_1365 <= _T_1364;
    _T_1366 <= _T_1365;
    _T_1367 <= _T_1366;
    _T_1368 <= _T_1367;
    _T_1369 <= _T_1368;
    _T_1370 <= _T_1369;
    _T_1371 <= _T_1370;
    _T_1372 <= _T_1371;
    _T_1373 <= _T_1372;
    _T_1374 <= _T_1373;
    _T_1375 <= _T_1374;
    _T_1376 <= _T_1375;
    _T_1377 <= _T_1376;
    _T_1378 <= _T_1377;
    _T_1379 <= _T_1378;
    _T_1380 <= _T_1379;
    _T_1381 <= _T_1380;
    _T_1382 <= _T_1381;
    _T_1383 <= _T_1382;
    _T_1384 <= _T_1383;
    _T_1385 <= _T_1384;
    _T_1386 <= _T_1385;
    _T_1387 <= _T_1386;
    _T_1388 <= _T_1387;
    _T_1389 <= _T_1388;
    _T_1390 <= _T_1389;
    _T_1391 <= _T_1390;
    _T_1392 <= _T_1391;
    _T_1393 <= _T_1392;
    _T_1394 <= _T_1393;
    _T_1395 <= _T_1394;
    _T_1396 <= _T_1395;
    _T_1397 <= _T_1396;
    _T_1398 <= _T_1397;
    _T_1399 <= _T_1398;
    _T_1400 <= _T_1399;
    _T_1401 <= _T_1400;
    _T_1402 <= _T_1401;
    _T_1403 <= _T_1402;
    _T_1404 <= _T_1403;
    _T_1405 <= _T_1404;
    _T_1406 <= _T_1405;
    _T_1407 <= _T_1406;
    _T_1408 <= _T_1407;
    _T_1409 <= _T_1408;
    _T_1410 <= _T_1409;
    _T_1411 <= _T_1410;
    _T_1412 <= _T_1411;
    _T_1413 <= _T_1412;
    _T_1414 <= _T_1413;
    _T_1415 <= _T_1414;
    _T_1416 <= _T_1415;
    _T_1417 <= _T_1416;
    _T_1418 <= _T_1417;
    _T_1419 <= _T_1418;
    _T_1420 <= _T_1419;
    _T_1421 <= _T_1420;
    _T_1422 <= _T_1421;
    _T_1423 <= _T_1422;
    _T_1424 <= _T_1423;
    _T_1425 <= _T_1424;
    _T_1426 <= _T_1425;
    _T_1427 <= _T_1426;
    _T_1428 <= _T_1427;
    _T_1429 <= _T_1428;
    _T_1430 <= _T_1429;
    _T_1431 <= _T_1430;
    _T_1432 <= _T_1431;
    _T_1433 <= _T_1432;
    _T_1434 <= _T_1433;
    _T_1435 <= _T_1434;
    _T_1436 <= _T_1435;
    _T_1437 <= _T_1436;
    _T_1438 <= _T_1437;
    _T_1439 <= _T_1438;
    _T_1440 <= _T_1439;
    _T_1441 <= _T_1440;
    _T_1442 <= _T_1441;
    _T_1443 <= _T_1442;
    _T_1444 <= _T_1443;
    _T_1445 <= _T_1444;
    _T_1446 <= _T_1445;
    _T_1447 <= _T_1446;
    _T_1448 <= _T_1447;
    _T_1449 <= _T_1448;
    _T_1450 <= _T_1449;
    _T_1451 <= _T_1450;
    _T_1452 <= _T_1451;
    _T_1453 <= _T_1452;
    _T_1454 <= _T_1453;
    _T_1455 <= _T_1454;
    _T_1456 <= _T_1455;
    _T_1457 <= _T_1456;
    _T_1458 <= _T_1457;
    _T_1459 <= _T_1458;
    _T_1460 <= _T_1459;
  end
endmodule
