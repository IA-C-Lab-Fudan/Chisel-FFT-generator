module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T; // @[Butterfly.scala 57:28]
  wire [63:0] _T_1; // @[Butterfly.scala 57:52]
  wire [63:0] _T_4; // @[Butterfly.scala 57:40]
  wire [63:0] _T_5; // @[Butterfly.scala 58:28]
  wire [63:0] _T_6; // @[Butterfly.scala 58:52]
  wire [63:0] _T_9; // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2; // @[Butterfly.scala 58:15]
  assign _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  assign _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  assign _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  assign _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  assign _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  assign _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  assign _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT128(
    input clk_in1_p,
    input clk_in1_n,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
    wire clock;
    clk_wiz_0 clk_wiz_0_inst0
       (
        // Clock out ports
        .clk_out1(clock),     // output clk_out1
       // Clock in ports
        .clk_in1_p(clk_in1_p),    // input clk_in1_p
        .clk_in1_n(clk_in1_n));    // input clk_in1_n
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [6:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [6:0] _T_1; // @[FFT.scala 42:16]
  wire [31:0] _GEN_2; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6; // @[FFT.scala 34:12]
  wire [31:0] _GEN_7; // @[FFT.scala 34:12]
  wire [31:0] _GEN_8; // @[FFT.scala 34:12]
  wire [31:0] _GEN_9; // @[FFT.scala 34:12]
  wire [31:0] _GEN_10; // @[FFT.scala 34:12]
  wire [31:0] _GEN_11; // @[FFT.scala 34:12]
  wire [31:0] _GEN_12; // @[FFT.scala 34:12]
  wire [31:0] _GEN_13; // @[FFT.scala 34:12]
  wire [31:0] _GEN_14; // @[FFT.scala 34:12]
  wire [31:0] _GEN_15; // @[FFT.scala 34:12]
  wire [31:0] _GEN_16; // @[FFT.scala 34:12]
  wire [31:0] _GEN_17; // @[FFT.scala 34:12]
  wire [31:0] _GEN_18; // @[FFT.scala 34:12]
  wire [31:0] _GEN_19; // @[FFT.scala 34:12]
  wire [31:0] _GEN_20; // @[FFT.scala 34:12]
  wire [31:0] _GEN_21; // @[FFT.scala 34:12]
  wire [31:0] _GEN_22; // @[FFT.scala 34:12]
  wire [31:0] _GEN_23; // @[FFT.scala 34:12]
  wire [31:0] _GEN_24; // @[FFT.scala 34:12]
  wire [31:0] _GEN_25; // @[FFT.scala 34:12]
  wire [31:0] _GEN_26; // @[FFT.scala 34:12]
  wire [31:0] _GEN_27; // @[FFT.scala 34:12]
  wire [31:0] _GEN_28; // @[FFT.scala 34:12]
  wire [31:0] _GEN_29; // @[FFT.scala 34:12]
  wire [31:0] _GEN_30; // @[FFT.scala 34:12]
  wire [31:0] _GEN_31; // @[FFT.scala 34:12]
  wire [31:0] _GEN_32; // @[FFT.scala 34:12]
  wire [31:0] _GEN_33; // @[FFT.scala 34:12]
  wire [31:0] _GEN_34; // @[FFT.scala 34:12]
  wire [31:0] _GEN_35; // @[FFT.scala 34:12]
  wire [31:0] _GEN_36; // @[FFT.scala 34:12]
  wire [31:0] _GEN_37; // @[FFT.scala 34:12]
  wire [31:0] _GEN_38; // @[FFT.scala 34:12]
  wire [31:0] _GEN_39; // @[FFT.scala 34:12]
  wire [31:0] _GEN_40; // @[FFT.scala 34:12]
  wire [31:0] _GEN_41; // @[FFT.scala 34:12]
  wire [31:0] _GEN_42; // @[FFT.scala 34:12]
  wire [31:0] _GEN_43; // @[FFT.scala 34:12]
  wire [31:0] _GEN_44; // @[FFT.scala 34:12]
  wire [31:0] _GEN_45; // @[FFT.scala 34:12]
  wire [31:0] _GEN_46; // @[FFT.scala 34:12]
  wire [31:0] _GEN_47; // @[FFT.scala 34:12]
  wire [31:0] _GEN_48; // @[FFT.scala 34:12]
  wire [31:0] _GEN_49; // @[FFT.scala 34:12]
  wire [31:0] _GEN_50; // @[FFT.scala 34:12]
  wire [31:0] _GEN_51; // @[FFT.scala 34:12]
  wire [31:0] _GEN_52; // @[FFT.scala 34:12]
  wire [31:0] _GEN_53; // @[FFT.scala 34:12]
  wire [31:0] _GEN_54; // @[FFT.scala 34:12]
  wire [31:0] _GEN_55; // @[FFT.scala 34:12]
  wire [31:0] _GEN_56; // @[FFT.scala 34:12]
  wire [31:0] _GEN_57; // @[FFT.scala 34:12]
  wire [31:0] _GEN_58; // @[FFT.scala 34:12]
  wire [31:0] _GEN_59; // @[FFT.scala 34:12]
  wire [31:0] _GEN_60; // @[FFT.scala 34:12]
  wire [31:0] _GEN_61; // @[FFT.scala 34:12]
  wire [31:0] _GEN_62; // @[FFT.scala 34:12]
  wire [31:0] _GEN_63; // @[FFT.scala 34:12]
  wire [31:0] _GEN_66; // @[FFT.scala 35:12]
  wire [31:0] _GEN_67; // @[FFT.scala 35:12]
  wire [31:0] _GEN_68; // @[FFT.scala 35:12]
  wire [31:0] _GEN_69; // @[FFT.scala 35:12]
  wire [31:0] _GEN_70; // @[FFT.scala 35:12]
  wire [31:0] _GEN_71; // @[FFT.scala 35:12]
  wire [31:0] _GEN_72; // @[FFT.scala 35:12]
  wire [31:0] _GEN_73; // @[FFT.scala 35:12]
  wire [31:0] _GEN_74; // @[FFT.scala 35:12]
  wire [31:0] _GEN_75; // @[FFT.scala 35:12]
  wire [31:0] _GEN_76; // @[FFT.scala 35:12]
  wire [31:0] _GEN_77; // @[FFT.scala 35:12]
  wire [31:0] _GEN_78; // @[FFT.scala 35:12]
  wire [31:0] _GEN_79; // @[FFT.scala 35:12]
  wire [31:0] _GEN_80; // @[FFT.scala 35:12]
  wire [31:0] _GEN_81; // @[FFT.scala 35:12]
  wire [31:0] _GEN_82; // @[FFT.scala 35:12]
  wire [31:0] _GEN_83; // @[FFT.scala 35:12]
  wire [31:0] _GEN_84; // @[FFT.scala 35:12]
  wire [31:0] _GEN_85; // @[FFT.scala 35:12]
  wire [31:0] _GEN_86; // @[FFT.scala 35:12]
  wire [31:0] _GEN_87; // @[FFT.scala 35:12]
  wire [31:0] _GEN_88; // @[FFT.scala 35:12]
  wire [31:0] _GEN_89; // @[FFT.scala 35:12]
  wire [31:0] _GEN_90; // @[FFT.scala 35:12]
  wire [31:0] _GEN_91; // @[FFT.scala 35:12]
  wire [31:0] _GEN_92; // @[FFT.scala 35:12]
  wire [31:0] _GEN_93; // @[FFT.scala 35:12]
  wire [31:0] _GEN_94; // @[FFT.scala 35:12]
  wire [31:0] _GEN_95; // @[FFT.scala 35:12]
  wire [31:0] _GEN_96; // @[FFT.scala 35:12]
  wire [31:0] _GEN_97; // @[FFT.scala 35:12]
  wire [31:0] _GEN_98; // @[FFT.scala 35:12]
  wire [31:0] _GEN_99; // @[FFT.scala 35:12]
  wire [31:0] _GEN_100; // @[FFT.scala 35:12]
  wire [31:0] _GEN_101; // @[FFT.scala 35:12]
  wire [31:0] _GEN_102; // @[FFT.scala 35:12]
  wire [31:0] _GEN_103; // @[FFT.scala 35:12]
  wire [31:0] _GEN_104; // @[FFT.scala 35:12]
  wire [31:0] _GEN_105; // @[FFT.scala 35:12]
  wire [31:0] _GEN_106; // @[FFT.scala 35:12]
  wire [31:0] _GEN_107; // @[FFT.scala 35:12]
  wire [31:0] _GEN_108; // @[FFT.scala 35:12]
  wire [31:0] _GEN_109; // @[FFT.scala 35:12]
  wire [31:0] _GEN_110; // @[FFT.scala 35:12]
  wire [31:0] _GEN_111; // @[FFT.scala 35:12]
  wire [31:0] _GEN_112; // @[FFT.scala 35:12]
  wire [31:0] _GEN_113; // @[FFT.scala 35:12]
  wire [31:0] _GEN_114; // @[FFT.scala 35:12]
  wire [31:0] _GEN_115; // @[FFT.scala 35:12]
  wire [31:0] _GEN_116; // @[FFT.scala 35:12]
  wire [31:0] _GEN_117; // @[FFT.scala 35:12]
  wire [31:0] _GEN_118; // @[FFT.scala 35:12]
  wire [31:0] _GEN_119; // @[FFT.scala 35:12]
  wire [31:0] _GEN_120; // @[FFT.scala 35:12]
  wire [31:0] _GEN_121; // @[FFT.scala 35:12]
  wire [31:0] _GEN_122; // @[FFT.scala 35:12]
  wire [31:0] _GEN_123; // @[FFT.scala 35:12]
  wire [31:0] _GEN_124; // @[FFT.scala 35:12]
  wire [31:0] _GEN_125; // @[FFT.scala 35:12]
  wire [31:0] _GEN_126; // @[FFT.scala 35:12]
  wire [31:0] _GEN_127; // @[FFT.scala 35:12]
  reg [31:0] _T_118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [31:0] _T_118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [31:0] _T_119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [31:0] _T_119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [31:0] _T_120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [31:0] _T_121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  wire [31:0] _GEN_322; // @[FFT.scala 34:12]
  wire [31:0] _GEN_323; // @[FFT.scala 34:12]
  wire [31:0] _GEN_324; // @[FFT.scala 34:12]
  wire [31:0] _GEN_325; // @[FFT.scala 34:12]
  wire [31:0] _GEN_326; // @[FFT.scala 34:12]
  wire [31:0] _GEN_327; // @[FFT.scala 34:12]
  wire [31:0] _GEN_328; // @[FFT.scala 34:12]
  wire [31:0] _GEN_329; // @[FFT.scala 34:12]
  wire [31:0] _GEN_330; // @[FFT.scala 34:12]
  wire [31:0] _GEN_331; // @[FFT.scala 34:12]
  wire [31:0] _GEN_332; // @[FFT.scala 34:12]
  wire [31:0] _GEN_333; // @[FFT.scala 34:12]
  wire [31:0] _GEN_334; // @[FFT.scala 34:12]
  wire [31:0] _GEN_335; // @[FFT.scala 34:12]
  wire [31:0] _GEN_336; // @[FFT.scala 34:12]
  wire [31:0] _GEN_337; // @[FFT.scala 34:12]
  wire [31:0] _GEN_338; // @[FFT.scala 34:12]
  wire [31:0] _GEN_339; // @[FFT.scala 34:12]
  wire [31:0] _GEN_340; // @[FFT.scala 34:12]
  wire [31:0] _GEN_341; // @[FFT.scala 34:12]
  wire [31:0] _GEN_342; // @[FFT.scala 34:12]
  wire [31:0] _GEN_343; // @[FFT.scala 34:12]
  wire [31:0] _GEN_344; // @[FFT.scala 34:12]
  wire [31:0] _GEN_345; // @[FFT.scala 34:12]
  wire [31:0] _GEN_346; // @[FFT.scala 34:12]
  wire [31:0] _GEN_347; // @[FFT.scala 34:12]
  wire [31:0] _GEN_348; // @[FFT.scala 34:12]
  wire [31:0] _GEN_349; // @[FFT.scala 34:12]
  wire [31:0] _GEN_350; // @[FFT.scala 34:12]
  wire [31:0] _GEN_351; // @[FFT.scala 34:12]
  wire [31:0] _GEN_354; // @[FFT.scala 35:12]
  wire [31:0] _GEN_355; // @[FFT.scala 35:12]
  wire [31:0] _GEN_356; // @[FFT.scala 35:12]
  wire [31:0] _GEN_357; // @[FFT.scala 35:12]
  wire [31:0] _GEN_358; // @[FFT.scala 35:12]
  wire [31:0] _GEN_359; // @[FFT.scala 35:12]
  wire [31:0] _GEN_360; // @[FFT.scala 35:12]
  wire [31:0] _GEN_361; // @[FFT.scala 35:12]
  wire [31:0] _GEN_362; // @[FFT.scala 35:12]
  wire [31:0] _GEN_363; // @[FFT.scala 35:12]
  wire [31:0] _GEN_364; // @[FFT.scala 35:12]
  wire [31:0] _GEN_365; // @[FFT.scala 35:12]
  wire [31:0] _GEN_366; // @[FFT.scala 35:12]
  wire [31:0] _GEN_367; // @[FFT.scala 35:12]
  wire [31:0] _GEN_368; // @[FFT.scala 35:12]
  wire [31:0] _GEN_369; // @[FFT.scala 35:12]
  wire [31:0] _GEN_370; // @[FFT.scala 35:12]
  wire [31:0] _GEN_371; // @[FFT.scala 35:12]
  wire [31:0] _GEN_372; // @[FFT.scala 35:12]
  wire [31:0] _GEN_373; // @[FFT.scala 35:12]
  wire [31:0] _GEN_374; // @[FFT.scala 35:12]
  wire [31:0] _GEN_375; // @[FFT.scala 35:12]
  wire [31:0] _GEN_376; // @[FFT.scala 35:12]
  wire [31:0] _GEN_377; // @[FFT.scala 35:12]
  wire [31:0] _GEN_378; // @[FFT.scala 35:12]
  wire [31:0] _GEN_379; // @[FFT.scala 35:12]
  wire [31:0] _GEN_380; // @[FFT.scala 35:12]
  wire [31:0] _GEN_381; // @[FFT.scala 35:12]
  wire [31:0] _GEN_382; // @[FFT.scala 35:12]
  wire [31:0] _GEN_383; // @[FFT.scala 35:12]
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  wire [31:0] _GEN_482; // @[FFT.scala 34:12]
  wire [31:0] _GEN_483; // @[FFT.scala 34:12]
  wire [31:0] _GEN_484; // @[FFT.scala 34:12]
  wire [31:0] _GEN_485; // @[FFT.scala 34:12]
  wire [31:0] _GEN_486; // @[FFT.scala 34:12]
  wire [31:0] _GEN_487; // @[FFT.scala 34:12]
  wire [31:0] _GEN_488; // @[FFT.scala 34:12]
  wire [31:0] _GEN_489; // @[FFT.scala 34:12]
  wire [31:0] _GEN_490; // @[FFT.scala 34:12]
  wire [31:0] _GEN_491; // @[FFT.scala 34:12]
  wire [31:0] _GEN_492; // @[FFT.scala 34:12]
  wire [31:0] _GEN_493; // @[FFT.scala 34:12]
  wire [31:0] _GEN_494; // @[FFT.scala 34:12]
  wire [31:0] _GEN_495; // @[FFT.scala 34:12]
  wire [31:0] _GEN_498; // @[FFT.scala 35:12]
  wire [31:0] _GEN_499; // @[FFT.scala 35:12]
  wire [31:0] _GEN_500; // @[FFT.scala 35:12]
  wire [31:0] _GEN_501; // @[FFT.scala 35:12]
  wire [31:0] _GEN_502; // @[FFT.scala 35:12]
  wire [31:0] _GEN_503; // @[FFT.scala 35:12]
  wire [31:0] _GEN_504; // @[FFT.scala 35:12]
  wire [31:0] _GEN_505; // @[FFT.scala 35:12]
  wire [31:0] _GEN_506; // @[FFT.scala 35:12]
  wire [31:0] _GEN_507; // @[FFT.scala 35:12]
  wire [31:0] _GEN_508; // @[FFT.scala 35:12]
  wire [31:0] _GEN_509; // @[FFT.scala 35:12]
  wire [31:0] _GEN_510; // @[FFT.scala 35:12]
  wire [31:0] _GEN_511; // @[FFT.scala 35:12]
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  wire [31:0] _GEN_562; // @[FFT.scala 34:12]
  wire [31:0] _GEN_563; // @[FFT.scala 34:12]
  wire [31:0] _GEN_564; // @[FFT.scala 34:12]
  wire [31:0] _GEN_565; // @[FFT.scala 34:12]
  wire [31:0] _GEN_566; // @[FFT.scala 34:12]
  wire [31:0] _GEN_567; // @[FFT.scala 34:12]
  wire [31:0] _GEN_570; // @[FFT.scala 35:12]
  wire [31:0] _GEN_571; // @[FFT.scala 35:12]
  wire [31:0] _GEN_572; // @[FFT.scala 35:12]
  wire [31:0] _GEN_573; // @[FFT.scala 35:12]
  wire [31:0] _GEN_574; // @[FFT.scala 35:12]
  wire [31:0] _GEN_575; // @[FFT.scala 35:12]
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  wire [31:0] _GEN_602; // @[FFT.scala 34:12]
  wire [31:0] _GEN_603; // @[FFT.scala 34:12]
  wire [31:0] _GEN_606; // @[FFT.scala 35:12]
  wire [31:0] _GEN_607; // @[FFT.scala 35:12]
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] out1D1_re; // @[FFT.scala 58:23]
  reg [31:0] _RAND_379;
  reg [31:0] out1D1_im; // @[FFT.scala 58:23]
  reg [31:0] _RAND_380;
  reg [31:0] _T_333_re; // @[FFT.scala 62:22]
  reg [31:0] _RAND_381;
  reg [31:0] _T_333_im; // @[FFT.scala 62:22]
  reg [31:0] _RAND_382;
  reg [31:0] _T_334_re; // @[FFT.scala 63:22]
  reg [31:0] _RAND_383;
  reg [31:0] _T_334_im; // @[FFT.scala 63:22]
  reg [31:0] _RAND_384;
  reg  _T_335; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg  _T_336; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg  _T_337; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg  _T_338; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg  _T_339; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg  _T_340; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg  _T_341; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg  _T_342; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg  _T_343; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg  _T_344; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg  _T_345; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg  _T_346; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg  _T_347; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg  _T_348; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg  _T_349; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg  _T_350; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg  _T_351; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg  _T_352; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg  _T_353; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg  _T_354; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg  _T_355; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg  _T_356; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg  _T_357; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg  _T_358; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg  _T_359; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg  _T_360; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg  _T_361; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg  _T_362; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg  _T_363; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg  _T_364; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg  _T_365; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg  _T_366; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg  _T_367; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg  _T_368; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg  _T_369; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg  _T_370; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg  _T_371; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg  _T_372; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg  _T_373; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg  _T_374; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg  _T_375; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg  _T_376; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg  _T_377; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg  _T_378; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg  _T_379; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg  _T_380; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg  _T_381; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg  _T_382; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg  _T_383; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg  _T_384; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg  _T_385; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg  _T_386; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg  _T_387; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg  _T_388; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg  _T_389; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg  _T_390; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg  _T_391; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg  _T_392; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg  _T_393; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg  _T_394; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg  _T_395; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg  _T_396; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg  _T_397; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg  _T_398; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg  _T_399; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg  _T_400; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg  _T_401; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg  _T_402; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg  _T_403; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg  _T_404; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg  _T_405; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg  _T_406; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg  _T_407; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg  _T_408; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg  _T_409; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg  _T_410; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg  _T_411; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg  _T_412; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg  _T_413; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg  _T_414; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg  _T_415; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg  _T_416; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg  _T_417; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg  _T_418; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg  _T_419; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg  _T_420; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg  _T_421; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg  _T_422; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg  _T_423; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg  _T_424; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg  _T_425; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg  _T_426; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg  _T_427; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg  _T_428; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg  _T_429; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg  _T_430; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg  _T_431; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg  _T_432; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg  _T_433; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg  _T_434; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg  _T_435; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg  _T_436; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg  _T_437; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg  _T_438; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg  _T_439; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg  _T_440; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg  _T_441; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg  _T_442; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg  _T_443; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg  _T_444; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg  _T_445; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg  _T_446; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg  _T_447; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg  _T_448; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg  _T_449; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg  _T_450; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg  _T_451; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg  _T_452; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg  _T_453; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg  _T_454; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg  _T_455; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg  _T_456; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg  _T_457; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg  _T_458; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg  _T_459; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg  _T_460; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg  _T_461; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg  _T_462; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign _T_1 = cnt + 7'h1; // @[FFT.scala 42:16]
  assign _GEN_2 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_3 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_2); // @[FFT.scala 34:12]
  assign _GEN_4 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_3); // @[FFT.scala 34:12]
  assign _GEN_5 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_4); // @[FFT.scala 34:12]
  assign _GEN_6 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_5); // @[FFT.scala 34:12]
  assign _GEN_7 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_6); // @[FFT.scala 34:12]
  assign _GEN_8 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_7); // @[FFT.scala 34:12]
  assign _GEN_9 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_8); // @[FFT.scala 34:12]
  assign _GEN_10 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_9); // @[FFT.scala 34:12]
  assign _GEN_11 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_10); // @[FFT.scala 34:12]
  assign _GEN_12 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_11); // @[FFT.scala 34:12]
  assign _GEN_13 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_12); // @[FFT.scala 34:12]
  assign _GEN_14 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_13); // @[FFT.scala 34:12]
  assign _GEN_15 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_14); // @[FFT.scala 34:12]
  assign _GEN_16 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_15); // @[FFT.scala 34:12]
  assign _GEN_17 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_16); // @[FFT.scala 34:12]
  assign _GEN_18 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_17); // @[FFT.scala 34:12]
  assign _GEN_19 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_18); // @[FFT.scala 34:12]
  assign _GEN_20 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_19); // @[FFT.scala 34:12]
  assign _GEN_21 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_20); // @[FFT.scala 34:12]
  assign _GEN_22 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_21); // @[FFT.scala 34:12]
  assign _GEN_23 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_22); // @[FFT.scala 34:12]
  assign _GEN_24 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_23); // @[FFT.scala 34:12]
  assign _GEN_25 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_24); // @[FFT.scala 34:12]
  assign _GEN_26 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_25); // @[FFT.scala 34:12]
  assign _GEN_27 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_26); // @[FFT.scala 34:12]
  assign _GEN_28 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_27); // @[FFT.scala 34:12]
  assign _GEN_29 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_28); // @[FFT.scala 34:12]
  assign _GEN_30 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_29); // @[FFT.scala 34:12]
  assign _GEN_31 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_30); // @[FFT.scala 34:12]
  assign _GEN_32 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_31); // @[FFT.scala 34:12]
  assign _GEN_33 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_32); // @[FFT.scala 34:12]
  assign _GEN_34 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_33); // @[FFT.scala 34:12]
  assign _GEN_35 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_34); // @[FFT.scala 34:12]
  assign _GEN_36 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_35); // @[FFT.scala 34:12]
  assign _GEN_37 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_36); // @[FFT.scala 34:12]
  assign _GEN_38 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_37); // @[FFT.scala 34:12]
  assign _GEN_39 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_38); // @[FFT.scala 34:12]
  assign _GEN_40 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_39); // @[FFT.scala 34:12]
  assign _GEN_41 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_40); // @[FFT.scala 34:12]
  assign _GEN_42 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_41); // @[FFT.scala 34:12]
  assign _GEN_43 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_42); // @[FFT.scala 34:12]
  assign _GEN_44 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_43); // @[FFT.scala 34:12]
  assign _GEN_45 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_44); // @[FFT.scala 34:12]
  assign _GEN_46 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_45); // @[FFT.scala 34:12]
  assign _GEN_47 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_46); // @[FFT.scala 34:12]
  assign _GEN_48 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_47); // @[FFT.scala 34:12]
  assign _GEN_49 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_48); // @[FFT.scala 34:12]
  assign _GEN_50 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_49); // @[FFT.scala 34:12]
  assign _GEN_51 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_50); // @[FFT.scala 34:12]
  assign _GEN_52 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_51); // @[FFT.scala 34:12]
  assign _GEN_53 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_52); // @[FFT.scala 34:12]
  assign _GEN_54 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_53); // @[FFT.scala 34:12]
  assign _GEN_55 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_54); // @[FFT.scala 34:12]
  assign _GEN_56 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_55); // @[FFT.scala 34:12]
  assign _GEN_57 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_56); // @[FFT.scala 34:12]
  assign _GEN_58 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_57); // @[FFT.scala 34:12]
  assign _GEN_59 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_58); // @[FFT.scala 34:12]
  assign _GEN_60 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_59); // @[FFT.scala 34:12]
  assign _GEN_61 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_60); // @[FFT.scala 34:12]
  assign _GEN_62 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_61); // @[FFT.scala 34:12]
  assign _GEN_63 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_62); // @[FFT.scala 34:12]
  assign _GEN_66 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_67 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_66); // @[FFT.scala 35:12]
  assign _GEN_68 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_67); // @[FFT.scala 35:12]
  assign _GEN_69 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_68); // @[FFT.scala 35:12]
  assign _GEN_70 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_69); // @[FFT.scala 35:12]
  assign _GEN_71 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_70); // @[FFT.scala 35:12]
  assign _GEN_72 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_71); // @[FFT.scala 35:12]
  assign _GEN_73 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_72); // @[FFT.scala 35:12]
  assign _GEN_74 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_73); // @[FFT.scala 35:12]
  assign _GEN_75 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_74); // @[FFT.scala 35:12]
  assign _GEN_76 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_75); // @[FFT.scala 35:12]
  assign _GEN_77 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_76); // @[FFT.scala 35:12]
  assign _GEN_78 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_77); // @[FFT.scala 35:12]
  assign _GEN_79 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_78); // @[FFT.scala 35:12]
  assign _GEN_80 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_79); // @[FFT.scala 35:12]
  assign _GEN_81 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_80); // @[FFT.scala 35:12]
  assign _GEN_82 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_81); // @[FFT.scala 35:12]
  assign _GEN_83 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_82); // @[FFT.scala 35:12]
  assign _GEN_84 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_83); // @[FFT.scala 35:12]
  assign _GEN_85 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_84); // @[FFT.scala 35:12]
  assign _GEN_86 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_85); // @[FFT.scala 35:12]
  assign _GEN_87 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_86); // @[FFT.scala 35:12]
  assign _GEN_88 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_87); // @[FFT.scala 35:12]
  assign _GEN_89 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_88); // @[FFT.scala 35:12]
  assign _GEN_90 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_89); // @[FFT.scala 35:12]
  assign _GEN_91 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_90); // @[FFT.scala 35:12]
  assign _GEN_92 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_91); // @[FFT.scala 35:12]
  assign _GEN_93 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_92); // @[FFT.scala 35:12]
  assign _GEN_94 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_93); // @[FFT.scala 35:12]
  assign _GEN_95 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_94); // @[FFT.scala 35:12]
  assign _GEN_96 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_95); // @[FFT.scala 35:12]
  assign _GEN_97 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_96); // @[FFT.scala 35:12]
  assign _GEN_98 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_97); // @[FFT.scala 35:12]
  assign _GEN_99 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_98); // @[FFT.scala 35:12]
  assign _GEN_100 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_99); // @[FFT.scala 35:12]
  assign _GEN_101 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_100); // @[FFT.scala 35:12]
  assign _GEN_102 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_101); // @[FFT.scala 35:12]
  assign _GEN_103 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_102); // @[FFT.scala 35:12]
  assign _GEN_104 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_103); // @[FFT.scala 35:12]
  assign _GEN_105 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_104); // @[FFT.scala 35:12]
  assign _GEN_106 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_105); // @[FFT.scala 35:12]
  assign _GEN_107 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_106); // @[FFT.scala 35:12]
  assign _GEN_108 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_107); // @[FFT.scala 35:12]
  assign _GEN_109 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_108); // @[FFT.scala 35:12]
  assign _GEN_110 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_109); // @[FFT.scala 35:12]
  assign _GEN_111 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_110); // @[FFT.scala 35:12]
  assign _GEN_112 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_111); // @[FFT.scala 35:12]
  assign _GEN_113 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_112); // @[FFT.scala 35:12]
  assign _GEN_114 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_113); // @[FFT.scala 35:12]
  assign _GEN_115 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_114); // @[FFT.scala 35:12]
  assign _GEN_116 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_115); // @[FFT.scala 35:12]
  assign _GEN_117 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_116); // @[FFT.scala 35:12]
  assign _GEN_118 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_117); // @[FFT.scala 35:12]
  assign _GEN_119 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_118); // @[FFT.scala 35:12]
  assign _GEN_120 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_119); // @[FFT.scala 35:12]
  assign _GEN_121 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_120); // @[FFT.scala 35:12]
  assign _GEN_122 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_121); // @[FFT.scala 35:12]
  assign _GEN_123 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_122); // @[FFT.scala 35:12]
  assign _GEN_124 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_123); // @[FFT.scala 35:12]
  assign _GEN_125 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_124); // @[FFT.scala 35:12]
  assign _GEN_126 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_125); // @[FFT.scala 35:12]
  assign _GEN_127 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_126); // @[FFT.scala 35:12]
  assign _GEN_322 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_323 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_322); // @[FFT.scala 34:12]
  assign _GEN_324 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_323); // @[FFT.scala 34:12]
  assign _GEN_325 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_324); // @[FFT.scala 34:12]
  assign _GEN_326 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_325); // @[FFT.scala 34:12]
  assign _GEN_327 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_326); // @[FFT.scala 34:12]
  assign _GEN_328 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_327); // @[FFT.scala 34:12]
  assign _GEN_329 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_328); // @[FFT.scala 34:12]
  assign _GEN_330 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_329); // @[FFT.scala 34:12]
  assign _GEN_331 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_330); // @[FFT.scala 34:12]
  assign _GEN_332 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_331); // @[FFT.scala 34:12]
  assign _GEN_333 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_332); // @[FFT.scala 34:12]
  assign _GEN_334 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_333); // @[FFT.scala 34:12]
  assign _GEN_335 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_334); // @[FFT.scala 34:12]
  assign _GEN_336 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_335); // @[FFT.scala 34:12]
  assign _GEN_337 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_336); // @[FFT.scala 34:12]
  assign _GEN_338 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_337); // @[FFT.scala 34:12]
  assign _GEN_339 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_338); // @[FFT.scala 34:12]
  assign _GEN_340 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_339); // @[FFT.scala 34:12]
  assign _GEN_341 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_340); // @[FFT.scala 34:12]
  assign _GEN_342 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_341); // @[FFT.scala 34:12]
  assign _GEN_343 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_342); // @[FFT.scala 34:12]
  assign _GEN_344 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_343); // @[FFT.scala 34:12]
  assign _GEN_345 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_344); // @[FFT.scala 34:12]
  assign _GEN_346 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_345); // @[FFT.scala 34:12]
  assign _GEN_347 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_346); // @[FFT.scala 34:12]
  assign _GEN_348 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_347); // @[FFT.scala 34:12]
  assign _GEN_349 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_348); // @[FFT.scala 34:12]
  assign _GEN_350 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_349); // @[FFT.scala 34:12]
  assign _GEN_351 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_350); // @[FFT.scala 34:12]
  assign _GEN_354 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_355 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_354); // @[FFT.scala 35:12]
  assign _GEN_356 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_355); // @[FFT.scala 35:12]
  assign _GEN_357 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_356); // @[FFT.scala 35:12]
  assign _GEN_358 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_357); // @[FFT.scala 35:12]
  assign _GEN_359 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_358); // @[FFT.scala 35:12]
  assign _GEN_360 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_359); // @[FFT.scala 35:12]
  assign _GEN_361 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_360); // @[FFT.scala 35:12]
  assign _GEN_362 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_361); // @[FFT.scala 35:12]
  assign _GEN_363 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_362); // @[FFT.scala 35:12]
  assign _GEN_364 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_363); // @[FFT.scala 35:12]
  assign _GEN_365 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_364); // @[FFT.scala 35:12]
  assign _GEN_366 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_365); // @[FFT.scala 35:12]
  assign _GEN_367 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_366); // @[FFT.scala 35:12]
  assign _GEN_368 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_367); // @[FFT.scala 35:12]
  assign _GEN_369 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_368); // @[FFT.scala 35:12]
  assign _GEN_370 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_369); // @[FFT.scala 35:12]
  assign _GEN_371 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_370); // @[FFT.scala 35:12]
  assign _GEN_372 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_371); // @[FFT.scala 35:12]
  assign _GEN_373 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_372); // @[FFT.scala 35:12]
  assign _GEN_374 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_373); // @[FFT.scala 35:12]
  assign _GEN_375 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_374); // @[FFT.scala 35:12]
  assign _GEN_376 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_375); // @[FFT.scala 35:12]
  assign _GEN_377 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_376); // @[FFT.scala 35:12]
  assign _GEN_378 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_377); // @[FFT.scala 35:12]
  assign _GEN_379 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_378); // @[FFT.scala 35:12]
  assign _GEN_380 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_379); // @[FFT.scala 35:12]
  assign _GEN_381 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_380); // @[FFT.scala 35:12]
  assign _GEN_382 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_381); // @[FFT.scala 35:12]
  assign _GEN_383 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_382); // @[FFT.scala 35:12]
  assign _GEN_482 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_483 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_482); // @[FFT.scala 34:12]
  assign _GEN_484 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_483); // @[FFT.scala 34:12]
  assign _GEN_485 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_484); // @[FFT.scala 34:12]
  assign _GEN_486 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_485); // @[FFT.scala 34:12]
  assign _GEN_487 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_486); // @[FFT.scala 34:12]
  assign _GEN_488 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_487); // @[FFT.scala 34:12]
  assign _GEN_489 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_488); // @[FFT.scala 34:12]
  assign _GEN_490 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_489); // @[FFT.scala 34:12]
  assign _GEN_491 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_490); // @[FFT.scala 34:12]
  assign _GEN_492 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_491); // @[FFT.scala 34:12]
  assign _GEN_493 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_492); // @[FFT.scala 34:12]
  assign _GEN_494 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_493); // @[FFT.scala 34:12]
  assign _GEN_495 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_494); // @[FFT.scala 34:12]
  assign _GEN_498 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_499 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_498); // @[FFT.scala 35:12]
  assign _GEN_500 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_499); // @[FFT.scala 35:12]
  assign _GEN_501 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_500); // @[FFT.scala 35:12]
  assign _GEN_502 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_501); // @[FFT.scala 35:12]
  assign _GEN_503 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_502); // @[FFT.scala 35:12]
  assign _GEN_504 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_503); // @[FFT.scala 35:12]
  assign _GEN_505 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_504); // @[FFT.scala 35:12]
  assign _GEN_506 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_505); // @[FFT.scala 35:12]
  assign _GEN_507 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_506); // @[FFT.scala 35:12]
  assign _GEN_508 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_507); // @[FFT.scala 35:12]
  assign _GEN_509 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_508); // @[FFT.scala 35:12]
  assign _GEN_510 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_509); // @[FFT.scala 35:12]
  assign _GEN_511 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_510); // @[FFT.scala 35:12]
  assign _GEN_562 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_563 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_562); // @[FFT.scala 34:12]
  assign _GEN_564 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_563); // @[FFT.scala 34:12]
  assign _GEN_565 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_564); // @[FFT.scala 34:12]
  assign _GEN_566 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_565); // @[FFT.scala 34:12]
  assign _GEN_567 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_566); // @[FFT.scala 34:12]
  assign _GEN_570 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_571 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_570); // @[FFT.scala 35:12]
  assign _GEN_572 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_571); // @[FFT.scala 35:12]
  assign _GEN_573 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_572); // @[FFT.scala 35:12]
  assign _GEN_574 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_573); // @[FFT.scala 35:12]
  assign _GEN_575 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_574); // @[FFT.scala 35:12]
  assign _GEN_602 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_603 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_602); // @[FFT.scala 34:12]
  assign _GEN_606 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_607 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_606); // @[FFT.scala 35:12]
  assign io_dOut1_re = _T_333_re; // @[FFT.scala 62:12]
  assign io_dOut1_im = _T_333_im; // @[FFT.scala 62:12]
  assign io_dOut2_re = _T_334_re; // @[FFT.scala 63:12]
  assign io_dOut2_im = _T_334_im; // @[FFT.scala 63:12]
  assign io_dout_valid = _T_462; // @[FFT.scala 64:17]
  assign Butterfly_io_in1_re = _T_181_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_181_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = io_dIn_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_63); // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_127); // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_214_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_214_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cnt[5]; // @[Butterfly.scala 113:17]
  assign Butterfly_1_io_in1_re = _T_250_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_250_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_351); // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_383); // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_267_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_267_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cnt[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_2_io_in1_re = _T_287_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_287_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_495); // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_511); // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_296_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_296_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cnt[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_3_io_in1_re = _T_308_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_308_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_567); // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_575); // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_313_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_313_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cnt[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_321_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_321_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_603); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_607); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_324_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_324_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cnt[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_330_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_330_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_332_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_332_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cnt[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_5_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_5_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_5_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_5_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_118_re = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_118_im = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_119_re = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_119_im = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_120_re = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_120_im = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_121_re = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_121_im = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_122_re = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_122_im = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_123_re = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_123_im = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_124_re = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_124_im = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_125_re = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_125_im = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_126_re = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_126_im = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_127_re = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_127_im = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_128_re = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_128_im = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_129_re = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_129_im = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_130_re = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_130_im = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_131_re = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_131_im = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_132_re = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_132_im = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_133_re = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_133_im = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_134_re = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_134_im = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_135_re = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_135_im = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_136_re = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_136_im = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_137_re = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_137_im = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_138_re = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_138_im = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_139_re = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_139_im = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_140_re = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_140_im = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_141_re = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_141_im = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_142_re = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_142_im = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_143_re = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_143_im = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_144_re = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_144_im = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_145_re = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_145_im = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_146_re = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_146_im = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_147_re = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_147_im = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_148_re = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_148_im = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_149_re = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_149_im = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_150_re = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_150_im = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_151_re = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_151_im = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_152_re = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_152_im = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_153_re = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_153_im = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_154_re = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_154_im = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_155_re = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_155_im = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_156_re = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_156_im = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_157_re = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_157_im = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_158_re = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_158_im = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_159_re = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_159_im = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_160_re = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_160_im = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_161_re = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_161_im = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_162_re = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_162_im = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_163_re = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_163_im = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_164_re = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_164_im = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_165_re = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_165_im = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_166_re = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_166_im = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_167_re = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_167_im = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_168_re = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_168_im = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_169_re = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_169_im = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_170_re = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_170_im = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_171_re = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_171_im = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_172_re = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_172_im = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_173_re = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_173_im = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_174_re = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_174_im = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_175_re = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_175_im = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_176_re = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_176_im = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_177_re = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_177_im = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_178_re = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_178_im = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_179_re = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_179_im = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_180_re = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_180_im = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_181_re = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_181_im = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_183_re = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_183_im = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_184_re = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_184_im = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_185_re = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_185_im = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_186_re = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_186_im = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_187_re = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_187_im = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_188_re = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_188_im = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_189_re = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_189_im = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_190_re = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_190_im = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_191_re = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_191_im = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_192_re = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_192_im = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_193_re = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_193_im = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_194_re = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_194_im = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_195_re = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_195_im = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_196_re = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_196_im = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_197_re = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_197_im = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_198_re = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_198_im = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_199_re = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_199_im = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_200_re = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_200_im = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_201_re = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_201_im = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_202_re = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_202_im = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_203_re = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_203_im = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_204_re = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_204_im = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_205_re = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_205_im = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_206_re = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_206_im = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_207_re = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_207_im = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_208_re = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_208_im = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_209_re = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_209_im = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_210_re = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_210_im = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_211_re = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_211_im = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_212_re = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_212_im = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_213_re = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_213_im = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_214_re = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_214_im = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_219_re = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_219_im = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_220_re = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_220_im = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_221_re = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_221_im = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_222_re = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_222_im = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_223_re = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_223_im = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_224_re = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_224_im = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_225_re = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_225_im = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_226_re = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_226_im = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_227_re = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_227_im = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_228_re = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_228_im = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_229_re = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_229_im = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_230_re = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_230_im = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_231_re = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_231_im = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_232_re = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_232_im = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_233_re = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_233_im = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_234_re = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_234_im = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_235_re = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_235_im = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_236_re = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_236_im = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_237_re = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_237_im = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_238_re = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_238_im = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_239_re = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_239_im = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_240_re = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_240_im = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_241_re = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_241_im = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_242_re = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_242_im = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_243_re = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_243_im = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_244_re = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_244_im = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_245_re = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_245_im = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_246_re = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_246_im = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_247_re = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_247_im = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_248_re = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_248_im = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_249_re = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_249_im = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_250_re = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_250_im = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_252_re = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_252_im = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_253_re = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_253_im = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_254_re = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_254_im = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_255_re = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_255_im = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_256_re = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_256_im = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_257_re = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_257_im = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_258_re = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_258_im = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_259_re = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_259_im = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_260_re = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_260_im = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_261_re = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_261_im = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_262_re = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_262_im = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_263_re = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_263_im = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_264_re = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_264_im = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_265_re = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_265_im = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_266_re = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_266_im = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_267_re = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_267_im = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_272_re = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_272_im = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_273_re = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_273_im = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_274_re = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_274_im = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_275_re = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_275_im = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_276_re = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_276_im = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_277_re = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_277_im = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_278_re = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_278_im = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_279_re = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_279_im = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_280_re = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_280_im = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_281_re = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_281_im = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_282_re = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_282_im = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_283_re = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_283_im = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_284_re = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_284_im = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_285_re = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_285_im = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_286_re = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_286_im = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_287_re = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_287_im = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_289_re = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_289_im = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_290_re = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_290_im = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_291_re = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_291_im = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_292_re = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_292_im = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_293_re = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_293_im = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_294_re = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_294_im = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_295_re = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_295_im = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_296_re = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_296_im = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_301_re = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_301_im = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_302_re = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_302_im = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_303_re = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_303_im = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_304_re = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_304_im = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_305_re = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_305_im = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_306_re = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_306_im = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_307_re = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_307_im = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_308_re = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_308_im = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_310_re = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_310_im = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_311_re = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_311_im = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_312_re = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_312_im = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_313_re = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_313_im = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_318_re = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_318_im = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_319_re = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_319_im = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_320_re = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_320_im = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_321_re = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_321_im = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_323_re = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_323_im = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_324_re = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_324_im = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_329_re = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_329_im = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_330_re = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_330_im = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_332_re = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_332_im = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  out1D1_re = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  out1D1_im = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_333_re = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_333_im = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_334_re = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_334_im = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_335 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_336 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_337 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_338 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_339 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_340 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_341 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_342 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_343 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_344 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_345 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_346 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_347 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_348 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_349 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_350 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_351 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_352 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_353 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_354 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_355 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_356 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_357 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_358 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_359 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_360 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_361 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_362 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_363 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_364 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_365 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_366 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_367 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_368 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_369 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_370 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_371 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_372 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_373 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_374 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_375 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_376 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_377 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_378 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_379 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_380 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_381 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_382 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_383 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_384 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_385 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_386 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_387 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_388 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_389 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_390 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_391 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_392 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_393 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_394 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_395 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_396 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_397 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_398 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_399 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_400 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_401 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_402 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_403 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_404 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_405 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_406 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_407 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_408 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_409 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_410 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_411 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_412 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_413 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_414 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_415 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_416 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_417 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_418 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_419 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_420 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_421 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_422 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_423 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_424 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_425 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_426 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_427 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_428 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_429 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_430 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_431 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_432 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_433 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_434 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_435 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_436 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_437 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_438 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_439 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_440 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_441 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_442 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_443 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_444 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_445 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_446 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_447 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_448 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_449 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_450 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_451 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_452 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_453 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_454 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_455 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_456 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_457 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_458 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_459 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_460 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_461 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_462 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 7'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    _T_118_re <= io_dIn_re;
    _T_118_im <= io_dIn_im;
    _T_119_re <= _T_118_re;
    _T_119_im <= _T_118_im;
    _T_120_re <= _T_119_re;
    _T_120_im <= _T_119_im;
    _T_121_re <= _T_120_re;
    _T_121_im <= _T_120_im;
    _T_122_re <= _T_121_re;
    _T_122_im <= _T_121_im;
    _T_123_re <= _T_122_re;
    _T_123_im <= _T_122_im;
    _T_124_re <= _T_123_re;
    _T_124_im <= _T_123_im;
    _T_125_re <= _T_124_re;
    _T_125_im <= _T_124_im;
    _T_126_re <= _T_125_re;
    _T_126_im <= _T_125_im;
    _T_127_re <= _T_126_re;
    _T_127_im <= _T_126_im;
    _T_128_re <= _T_127_re;
    _T_128_im <= _T_127_im;
    _T_129_re <= _T_128_re;
    _T_129_im <= _T_128_im;
    _T_130_re <= _T_129_re;
    _T_130_im <= _T_129_im;
    _T_131_re <= _T_130_re;
    _T_131_im <= _T_130_im;
    _T_132_re <= _T_131_re;
    _T_132_im <= _T_131_im;
    _T_133_re <= _T_132_re;
    _T_133_im <= _T_132_im;
    _T_134_re <= _T_133_re;
    _T_134_im <= _T_133_im;
    _T_135_re <= _T_134_re;
    _T_135_im <= _T_134_im;
    _T_136_re <= _T_135_re;
    _T_136_im <= _T_135_im;
    _T_137_re <= _T_136_re;
    _T_137_im <= _T_136_im;
    _T_138_re <= _T_137_re;
    _T_138_im <= _T_137_im;
    _T_139_re <= _T_138_re;
    _T_139_im <= _T_138_im;
    _T_140_re <= _T_139_re;
    _T_140_im <= _T_139_im;
    _T_141_re <= _T_140_re;
    _T_141_im <= _T_140_im;
    _T_142_re <= _T_141_re;
    _T_142_im <= _T_141_im;
    _T_143_re <= _T_142_re;
    _T_143_im <= _T_142_im;
    _T_144_re <= _T_143_re;
    _T_144_im <= _T_143_im;
    _T_145_re <= _T_144_re;
    _T_145_im <= _T_144_im;
    _T_146_re <= _T_145_re;
    _T_146_im <= _T_145_im;
    _T_147_re <= _T_146_re;
    _T_147_im <= _T_146_im;
    _T_148_re <= _T_147_re;
    _T_148_im <= _T_147_im;
    _T_149_re <= _T_148_re;
    _T_149_im <= _T_148_im;
    _T_150_re <= _T_149_re;
    _T_150_im <= _T_149_im;
    _T_151_re <= _T_150_re;
    _T_151_im <= _T_150_im;
    _T_152_re <= _T_151_re;
    _T_152_im <= _T_151_im;
    _T_153_re <= _T_152_re;
    _T_153_im <= _T_152_im;
    _T_154_re <= _T_153_re;
    _T_154_im <= _T_153_im;
    _T_155_re <= _T_154_re;
    _T_155_im <= _T_154_im;
    _T_156_re <= _T_155_re;
    _T_156_im <= _T_155_im;
    _T_157_re <= _T_156_re;
    _T_157_im <= _T_156_im;
    _T_158_re <= _T_157_re;
    _T_158_im <= _T_157_im;
    _T_159_re <= _T_158_re;
    _T_159_im <= _T_158_im;
    _T_160_re <= _T_159_re;
    _T_160_im <= _T_159_im;
    _T_161_re <= _T_160_re;
    _T_161_im <= _T_160_im;
    _T_162_re <= _T_161_re;
    _T_162_im <= _T_161_im;
    _T_163_re <= _T_162_re;
    _T_163_im <= _T_162_im;
    _T_164_re <= _T_163_re;
    _T_164_im <= _T_163_im;
    _T_165_re <= _T_164_re;
    _T_165_im <= _T_164_im;
    _T_166_re <= _T_165_re;
    _T_166_im <= _T_165_im;
    _T_167_re <= _T_166_re;
    _T_167_im <= _T_166_im;
    _T_168_re <= _T_167_re;
    _T_168_im <= _T_167_im;
    _T_169_re <= _T_168_re;
    _T_169_im <= _T_168_im;
    _T_170_re <= _T_169_re;
    _T_170_im <= _T_169_im;
    _T_171_re <= _T_170_re;
    _T_171_im <= _T_170_im;
    _T_172_re <= _T_171_re;
    _T_172_im <= _T_171_im;
    _T_173_re <= _T_172_re;
    _T_173_im <= _T_172_im;
    _T_174_re <= _T_173_re;
    _T_174_im <= _T_173_im;
    _T_175_re <= _T_174_re;
    _T_175_im <= _T_174_im;
    _T_176_re <= _T_175_re;
    _T_176_im <= _T_175_im;
    _T_177_re <= _T_176_re;
    _T_177_im <= _T_176_im;
    _T_178_re <= _T_177_re;
    _T_178_im <= _T_177_im;
    _T_179_re <= _T_178_re;
    _T_179_im <= _T_178_im;
    _T_180_re <= _T_179_re;
    _T_180_im <= _T_179_im;
    _T_181_re <= _T_180_re;
    _T_181_im <= _T_180_im;
    _T_183_re <= Butterfly_io_out2_re;
    _T_183_im <= Butterfly_io_out2_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_219_re <= Switch_io_out1_re;
    _T_219_im <= Switch_io_out1_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_252_re <= Butterfly_1_io_out2_re;
    _T_252_im <= Butterfly_1_io_out2_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_272_re <= Switch_1_io_out1_re;
    _T_272_im <= Switch_1_io_out1_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_289_re <= Butterfly_2_io_out2_re;
    _T_289_im <= Butterfly_2_io_out2_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_301_re <= Switch_2_io_out1_re;
    _T_301_im <= Switch_2_io_out1_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_310_re <= Butterfly_3_io_out2_re;
    _T_310_im <= Butterfly_3_io_out2_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_318_re <= Switch_3_io_out1_re;
    _T_318_im <= Switch_3_io_out1_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_323_re <= Butterfly_4_io_out2_re;
    _T_323_im <= Butterfly_4_io_out2_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_329_re <= Switch_4_io_out1_re;
    _T_329_im <= Switch_4_io_out1_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_332_re <= Butterfly_5_io_out2_re;
    _T_332_im <= Butterfly_5_io_out2_im;
    out1D1_re <= Switch_5_io_out1_re;
    out1D1_im <= Switch_5_io_out1_im;
    _T_333_re <= ComplexAdd_io_res_re;
    _T_333_im <= ComplexAdd_io_res_im;
    _T_334_re <= ComplexSub_io_res_re;
    _T_334_im <= ComplexSub_io_res_im;
    _T_335 <= io_din_valid;
    _T_336 <= _T_335;
    _T_337 <= _T_336;
    _T_338 <= _T_337;
    _T_339 <= _T_338;
    _T_340 <= _T_339;
    _T_341 <= _T_340;
    _T_342 <= _T_341;
    _T_343 <= _T_342;
    _T_344 <= _T_343;
    _T_345 <= _T_344;
    _T_346 <= _T_345;
    _T_347 <= _T_346;
    _T_348 <= _T_347;
    _T_349 <= _T_348;
    _T_350 <= _T_349;
    _T_351 <= _T_350;
    _T_352 <= _T_351;
    _T_353 <= _T_352;
    _T_354 <= _T_353;
    _T_355 <= _T_354;
    _T_356 <= _T_355;
    _T_357 <= _T_356;
    _T_358 <= _T_357;
    _T_359 <= _T_358;
    _T_360 <= _T_359;
    _T_361 <= _T_360;
    _T_362 <= _T_361;
    _T_363 <= _T_362;
    _T_364 <= _T_363;
    _T_365 <= _T_364;
    _T_366 <= _T_365;
    _T_367 <= _T_366;
    _T_368 <= _T_367;
    _T_369 <= _T_368;
    _T_370 <= _T_369;
    _T_371 <= _T_370;
    _T_372 <= _T_371;
    _T_373 <= _T_372;
    _T_374 <= _T_373;
    _T_375 <= _T_374;
    _T_376 <= _T_375;
    _T_377 <= _T_376;
    _T_378 <= _T_377;
    _T_379 <= _T_378;
    _T_380 <= _T_379;
    _T_381 <= _T_380;
    _T_382 <= _T_381;
    _T_383 <= _T_382;
    _T_384 <= _T_383;
    _T_385 <= _T_384;
    _T_386 <= _T_385;
    _T_387 <= _T_386;
    _T_388 <= _T_387;
    _T_389 <= _T_388;
    _T_390 <= _T_389;
    _T_391 <= _T_390;
    _T_392 <= _T_391;
    _T_393 <= _T_392;
    _T_394 <= _T_393;
    _T_395 <= _T_394;
    _T_396 <= _T_395;
    _T_397 <= _T_396;
    _T_398 <= _T_397;
    _T_399 <= _T_398;
    _T_400 <= _T_399;
    _T_401 <= _T_400;
    _T_402 <= _T_401;
    _T_403 <= _T_402;
    _T_404 <= _T_403;
    _T_405 <= _T_404;
    _T_406 <= _T_405;
    _T_407 <= _T_406;
    _T_408 <= _T_407;
    _T_409 <= _T_408;
    _T_410 <= _T_409;
    _T_411 <= _T_410;
    _T_412 <= _T_411;
    _T_413 <= _T_412;
    _T_414 <= _T_413;
    _T_415 <= _T_414;
    _T_416 <= _T_415;
    _T_417 <= _T_416;
    _T_418 <= _T_417;
    _T_419 <= _T_418;
    _T_420 <= _T_419;
    _T_421 <= _T_420;
    _T_422 <= _T_421;
    _T_423 <= _T_422;
    _T_424 <= _T_423;
    _T_425 <= _T_424;
    _T_426 <= _T_425;
    _T_427 <= _T_426;
    _T_428 <= _T_427;
    _T_429 <= _T_428;
    _T_430 <= _T_429;
    _T_431 <= _T_430;
    _T_432 <= _T_431;
    _T_433 <= _T_432;
    _T_434 <= _T_433;
    _T_435 <= _T_434;
    _T_436 <= _T_435;
    _T_437 <= _T_436;
    _T_438 <= _T_437;
    _T_439 <= _T_438;
    _T_440 <= _T_439;
    _T_441 <= _T_440;
    _T_442 <= _T_441;
    _T_443 <= _T_442;
    _T_444 <= _T_443;
    _T_445 <= _T_444;
    _T_446 <= _T_445;
    _T_447 <= _T_446;
    _T_448 <= _T_447;
    _T_449 <= _T_448;
    _T_450 <= _T_449;
    _T_451 <= _T_450;
    _T_452 <= _T_451;
    _T_453 <= _T_452;
    _T_454 <= _T_453;
    _T_455 <= _T_454;
    _T_456 <= _T_455;
    _T_457 <= _T_456;
    _T_458 <= _T_457;
    _T_459 <= _T_458;
    _T_460 <= _T_459;
    _T_461 <= _T_460;
    _T_462 <= _T_461;
  end
endmodule
