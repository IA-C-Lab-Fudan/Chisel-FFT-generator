module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T; // @[Butterfly.scala 57:28]
  wire [63:0] _T_1; // @[Butterfly.scala 57:52]
  wire [63:0] _T_4; // @[Butterfly.scala 57:40]
  wire [63:0] _T_5; // @[Butterfly.scala 58:28]
  wire [63:0] _T_6; // @[Butterfly.scala 58:52]
  wire [63:0] _T_9; // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2; // @[Butterfly.scala 58:15]
  assign _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  assign _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  assign _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  assign _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  assign _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  assign _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  assign _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT1024(
    input clk_in1_p,
    input clk_in1_n,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
    wire clock;
    clk_wiz_0 clk_wiz_0_inst0
       (
        // Clock out ports
        .clk_out1(clock),     // output clk_out1
       // Clock in ports
        .clk_in1_p(clk_in1_p),    // input clk_in1_p
        .clk_in1_n(clk_in1_n));    // input clk_in1_n
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_8_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_8_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_8_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [9:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [9:0] _T_1; // @[FFT.scala 42:16]
  reg [9:0] cntD1; // @[FFT.scala 44:22]
  reg [31:0] _RAND_1;
  wire [31:0] _GEN_2; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6; // @[FFT.scala 34:12]
  wire [31:0] _GEN_7; // @[FFT.scala 34:12]
  wire [31:0] _GEN_8; // @[FFT.scala 34:12]
  wire [31:0] _GEN_9; // @[FFT.scala 34:12]
  wire [31:0] _GEN_10; // @[FFT.scala 34:12]
  wire [31:0] _GEN_11; // @[FFT.scala 34:12]
  wire [31:0] _GEN_12; // @[FFT.scala 34:12]
  wire [31:0] _GEN_13; // @[FFT.scala 34:12]
  wire [31:0] _GEN_14; // @[FFT.scala 34:12]
  wire [31:0] _GEN_15; // @[FFT.scala 34:12]
  wire [31:0] _GEN_16; // @[FFT.scala 34:12]
  wire [31:0] _GEN_17; // @[FFT.scala 34:12]
  wire [31:0] _GEN_18; // @[FFT.scala 34:12]
  wire [31:0] _GEN_19; // @[FFT.scala 34:12]
  wire [31:0] _GEN_20; // @[FFT.scala 34:12]
  wire [31:0] _GEN_21; // @[FFT.scala 34:12]
  wire [31:0] _GEN_22; // @[FFT.scala 34:12]
  wire [31:0] _GEN_23; // @[FFT.scala 34:12]
  wire [31:0] _GEN_24; // @[FFT.scala 34:12]
  wire [31:0] _GEN_25; // @[FFT.scala 34:12]
  wire [31:0] _GEN_26; // @[FFT.scala 34:12]
  wire [31:0] _GEN_27; // @[FFT.scala 34:12]
  wire [31:0] _GEN_28; // @[FFT.scala 34:12]
  wire [31:0] _GEN_29; // @[FFT.scala 34:12]
  wire [31:0] _GEN_30; // @[FFT.scala 34:12]
  wire [31:0] _GEN_31; // @[FFT.scala 34:12]
  wire [31:0] _GEN_32; // @[FFT.scala 34:12]
  wire [31:0] _GEN_33; // @[FFT.scala 34:12]
  wire [31:0] _GEN_34; // @[FFT.scala 34:12]
  wire [31:0] _GEN_35; // @[FFT.scala 34:12]
  wire [31:0] _GEN_36; // @[FFT.scala 34:12]
  wire [31:0] _GEN_37; // @[FFT.scala 34:12]
  wire [31:0] _GEN_38; // @[FFT.scala 34:12]
  wire [31:0] _GEN_39; // @[FFT.scala 34:12]
  wire [31:0] _GEN_40; // @[FFT.scala 34:12]
  wire [31:0] _GEN_41; // @[FFT.scala 34:12]
  wire [31:0] _GEN_42; // @[FFT.scala 34:12]
  wire [31:0] _GEN_43; // @[FFT.scala 34:12]
  wire [31:0] _GEN_44; // @[FFT.scala 34:12]
  wire [31:0] _GEN_45; // @[FFT.scala 34:12]
  wire [31:0] _GEN_46; // @[FFT.scala 34:12]
  wire [31:0] _GEN_47; // @[FFT.scala 34:12]
  wire [31:0] _GEN_48; // @[FFT.scala 34:12]
  wire [31:0] _GEN_49; // @[FFT.scala 34:12]
  wire [31:0] _GEN_50; // @[FFT.scala 34:12]
  wire [31:0] _GEN_51; // @[FFT.scala 34:12]
  wire [31:0] _GEN_52; // @[FFT.scala 34:12]
  wire [31:0] _GEN_53; // @[FFT.scala 34:12]
  wire [31:0] _GEN_54; // @[FFT.scala 34:12]
  wire [31:0] _GEN_55; // @[FFT.scala 34:12]
  wire [31:0] _GEN_56; // @[FFT.scala 34:12]
  wire [31:0] _GEN_57; // @[FFT.scala 34:12]
  wire [31:0] _GEN_58; // @[FFT.scala 34:12]
  wire [31:0] _GEN_59; // @[FFT.scala 34:12]
  wire [31:0] _GEN_60; // @[FFT.scala 34:12]
  wire [31:0] _GEN_61; // @[FFT.scala 34:12]
  wire [31:0] _GEN_62; // @[FFT.scala 34:12]
  wire [31:0] _GEN_63; // @[FFT.scala 34:12]
  wire [31:0] _GEN_64; // @[FFT.scala 34:12]
  wire [31:0] _GEN_65; // @[FFT.scala 34:12]
  wire [31:0] _GEN_66; // @[FFT.scala 34:12]
  wire [31:0] _GEN_67; // @[FFT.scala 34:12]
  wire [31:0] _GEN_68; // @[FFT.scala 34:12]
  wire [31:0] _GEN_69; // @[FFT.scala 34:12]
  wire [31:0] _GEN_70; // @[FFT.scala 34:12]
  wire [31:0] _GEN_71; // @[FFT.scala 34:12]
  wire [31:0] _GEN_72; // @[FFT.scala 34:12]
  wire [31:0] _GEN_73; // @[FFT.scala 34:12]
  wire [31:0] _GEN_74; // @[FFT.scala 34:12]
  wire [31:0] _GEN_75; // @[FFT.scala 34:12]
  wire [31:0] _GEN_76; // @[FFT.scala 34:12]
  wire [31:0] _GEN_77; // @[FFT.scala 34:12]
  wire [31:0] _GEN_78; // @[FFT.scala 34:12]
  wire [31:0] _GEN_79; // @[FFT.scala 34:12]
  wire [31:0] _GEN_80; // @[FFT.scala 34:12]
  wire [31:0] _GEN_81; // @[FFT.scala 34:12]
  wire [31:0] _GEN_82; // @[FFT.scala 34:12]
  wire [31:0] _GEN_83; // @[FFT.scala 34:12]
  wire [31:0] _GEN_84; // @[FFT.scala 34:12]
  wire [31:0] _GEN_85; // @[FFT.scala 34:12]
  wire [31:0] _GEN_86; // @[FFT.scala 34:12]
  wire [31:0] _GEN_87; // @[FFT.scala 34:12]
  wire [31:0] _GEN_88; // @[FFT.scala 34:12]
  wire [31:0] _GEN_89; // @[FFT.scala 34:12]
  wire [31:0] _GEN_90; // @[FFT.scala 34:12]
  wire [31:0] _GEN_91; // @[FFT.scala 34:12]
  wire [31:0] _GEN_92; // @[FFT.scala 34:12]
  wire [31:0] _GEN_93; // @[FFT.scala 34:12]
  wire [31:0] _GEN_94; // @[FFT.scala 34:12]
  wire [31:0] _GEN_95; // @[FFT.scala 34:12]
  wire [31:0] _GEN_96; // @[FFT.scala 34:12]
  wire [31:0] _GEN_97; // @[FFT.scala 34:12]
  wire [31:0] _GEN_98; // @[FFT.scala 34:12]
  wire [31:0] _GEN_99; // @[FFT.scala 34:12]
  wire [31:0] _GEN_100; // @[FFT.scala 34:12]
  wire [31:0] _GEN_101; // @[FFT.scala 34:12]
  wire [31:0] _GEN_102; // @[FFT.scala 34:12]
  wire [31:0] _GEN_103; // @[FFT.scala 34:12]
  wire [31:0] _GEN_104; // @[FFT.scala 34:12]
  wire [31:0] _GEN_105; // @[FFT.scala 34:12]
  wire [31:0] _GEN_106; // @[FFT.scala 34:12]
  wire [31:0] _GEN_107; // @[FFT.scala 34:12]
  wire [31:0] _GEN_108; // @[FFT.scala 34:12]
  wire [31:0] _GEN_109; // @[FFT.scala 34:12]
  wire [31:0] _GEN_110; // @[FFT.scala 34:12]
  wire [31:0] _GEN_111; // @[FFT.scala 34:12]
  wire [31:0] _GEN_112; // @[FFT.scala 34:12]
  wire [31:0] _GEN_113; // @[FFT.scala 34:12]
  wire [31:0] _GEN_114; // @[FFT.scala 34:12]
  wire [31:0] _GEN_115; // @[FFT.scala 34:12]
  wire [31:0] _GEN_116; // @[FFT.scala 34:12]
  wire [31:0] _GEN_117; // @[FFT.scala 34:12]
  wire [31:0] _GEN_118; // @[FFT.scala 34:12]
  wire [31:0] _GEN_119; // @[FFT.scala 34:12]
  wire [31:0] _GEN_120; // @[FFT.scala 34:12]
  wire [31:0] _GEN_121; // @[FFT.scala 34:12]
  wire [31:0] _GEN_122; // @[FFT.scala 34:12]
  wire [31:0] _GEN_123; // @[FFT.scala 34:12]
  wire [31:0] _GEN_124; // @[FFT.scala 34:12]
  wire [31:0] _GEN_125; // @[FFT.scala 34:12]
  wire [31:0] _GEN_126; // @[FFT.scala 34:12]
  wire [31:0] _GEN_127; // @[FFT.scala 34:12]
  wire [31:0] _GEN_128; // @[FFT.scala 34:12]
  wire [31:0] _GEN_129; // @[FFT.scala 34:12]
  wire [31:0] _GEN_130; // @[FFT.scala 34:12]
  wire [31:0] _GEN_131; // @[FFT.scala 34:12]
  wire [31:0] _GEN_132; // @[FFT.scala 34:12]
  wire [31:0] _GEN_133; // @[FFT.scala 34:12]
  wire [31:0] _GEN_134; // @[FFT.scala 34:12]
  wire [31:0] _GEN_135; // @[FFT.scala 34:12]
  wire [31:0] _GEN_136; // @[FFT.scala 34:12]
  wire [31:0] _GEN_137; // @[FFT.scala 34:12]
  wire [31:0] _GEN_138; // @[FFT.scala 34:12]
  wire [31:0] _GEN_139; // @[FFT.scala 34:12]
  wire [31:0] _GEN_140; // @[FFT.scala 34:12]
  wire [31:0] _GEN_141; // @[FFT.scala 34:12]
  wire [31:0] _GEN_142; // @[FFT.scala 34:12]
  wire [31:0] _GEN_143; // @[FFT.scala 34:12]
  wire [31:0] _GEN_144; // @[FFT.scala 34:12]
  wire [31:0] _GEN_145; // @[FFT.scala 34:12]
  wire [31:0] _GEN_146; // @[FFT.scala 34:12]
  wire [31:0] _GEN_147; // @[FFT.scala 34:12]
  wire [31:0] _GEN_148; // @[FFT.scala 34:12]
  wire [31:0] _GEN_149; // @[FFT.scala 34:12]
  wire [31:0] _GEN_150; // @[FFT.scala 34:12]
  wire [31:0] _GEN_151; // @[FFT.scala 34:12]
  wire [31:0] _GEN_152; // @[FFT.scala 34:12]
  wire [31:0] _GEN_153; // @[FFT.scala 34:12]
  wire [31:0] _GEN_154; // @[FFT.scala 34:12]
  wire [31:0] _GEN_155; // @[FFT.scala 34:12]
  wire [31:0] _GEN_156; // @[FFT.scala 34:12]
  wire [31:0] _GEN_157; // @[FFT.scala 34:12]
  wire [31:0] _GEN_158; // @[FFT.scala 34:12]
  wire [31:0] _GEN_159; // @[FFT.scala 34:12]
  wire [31:0] _GEN_160; // @[FFT.scala 34:12]
  wire [31:0] _GEN_161; // @[FFT.scala 34:12]
  wire [31:0] _GEN_162; // @[FFT.scala 34:12]
  wire [31:0] _GEN_163; // @[FFT.scala 34:12]
  wire [31:0] _GEN_164; // @[FFT.scala 34:12]
  wire [31:0] _GEN_165; // @[FFT.scala 34:12]
  wire [31:0] _GEN_166; // @[FFT.scala 34:12]
  wire [31:0] _GEN_167; // @[FFT.scala 34:12]
  wire [31:0] _GEN_168; // @[FFT.scala 34:12]
  wire [31:0] _GEN_169; // @[FFT.scala 34:12]
  wire [31:0] _GEN_170; // @[FFT.scala 34:12]
  wire [31:0] _GEN_171; // @[FFT.scala 34:12]
  wire [31:0] _GEN_172; // @[FFT.scala 34:12]
  wire [31:0] _GEN_173; // @[FFT.scala 34:12]
  wire [31:0] _GEN_174; // @[FFT.scala 34:12]
  wire [31:0] _GEN_175; // @[FFT.scala 34:12]
  wire [31:0] _GEN_176; // @[FFT.scala 34:12]
  wire [31:0] _GEN_177; // @[FFT.scala 34:12]
  wire [31:0] _GEN_178; // @[FFT.scala 34:12]
  wire [31:0] _GEN_179; // @[FFT.scala 34:12]
  wire [31:0] _GEN_180; // @[FFT.scala 34:12]
  wire [31:0] _GEN_181; // @[FFT.scala 34:12]
  wire [31:0] _GEN_182; // @[FFT.scala 34:12]
  wire [31:0] _GEN_183; // @[FFT.scala 34:12]
  wire [31:0] _GEN_184; // @[FFT.scala 34:12]
  wire [31:0] _GEN_185; // @[FFT.scala 34:12]
  wire [31:0] _GEN_186; // @[FFT.scala 34:12]
  wire [31:0] _GEN_187; // @[FFT.scala 34:12]
  wire [31:0] _GEN_188; // @[FFT.scala 34:12]
  wire [31:0] _GEN_189; // @[FFT.scala 34:12]
  wire [31:0] _GEN_190; // @[FFT.scala 34:12]
  wire [31:0] _GEN_191; // @[FFT.scala 34:12]
  wire [31:0] _GEN_192; // @[FFT.scala 34:12]
  wire [31:0] _GEN_193; // @[FFT.scala 34:12]
  wire [31:0] _GEN_194; // @[FFT.scala 34:12]
  wire [31:0] _GEN_195; // @[FFT.scala 34:12]
  wire [31:0] _GEN_196; // @[FFT.scala 34:12]
  wire [31:0] _GEN_197; // @[FFT.scala 34:12]
  wire [31:0] _GEN_198; // @[FFT.scala 34:12]
  wire [31:0] _GEN_199; // @[FFT.scala 34:12]
  wire [31:0] _GEN_200; // @[FFT.scala 34:12]
  wire [31:0] _GEN_201; // @[FFT.scala 34:12]
  wire [31:0] _GEN_202; // @[FFT.scala 34:12]
  wire [31:0] _GEN_203; // @[FFT.scala 34:12]
  wire [31:0] _GEN_204; // @[FFT.scala 34:12]
  wire [31:0] _GEN_205; // @[FFT.scala 34:12]
  wire [31:0] _GEN_206; // @[FFT.scala 34:12]
  wire [31:0] _GEN_207; // @[FFT.scala 34:12]
  wire [31:0] _GEN_208; // @[FFT.scala 34:12]
  wire [31:0] _GEN_209; // @[FFT.scala 34:12]
  wire [31:0] _GEN_210; // @[FFT.scala 34:12]
  wire [31:0] _GEN_211; // @[FFT.scala 34:12]
  wire [31:0] _GEN_212; // @[FFT.scala 34:12]
  wire [31:0] _GEN_213; // @[FFT.scala 34:12]
  wire [31:0] _GEN_214; // @[FFT.scala 34:12]
  wire [31:0] _GEN_215; // @[FFT.scala 34:12]
  wire [31:0] _GEN_216; // @[FFT.scala 34:12]
  wire [31:0] _GEN_217; // @[FFT.scala 34:12]
  wire [31:0] _GEN_218; // @[FFT.scala 34:12]
  wire [31:0] _GEN_219; // @[FFT.scala 34:12]
  wire [31:0] _GEN_220; // @[FFT.scala 34:12]
  wire [31:0] _GEN_221; // @[FFT.scala 34:12]
  wire [31:0] _GEN_222; // @[FFT.scala 34:12]
  wire [31:0] _GEN_223; // @[FFT.scala 34:12]
  wire [31:0] _GEN_224; // @[FFT.scala 34:12]
  wire [31:0] _GEN_225; // @[FFT.scala 34:12]
  wire [31:0] _GEN_226; // @[FFT.scala 34:12]
  wire [31:0] _GEN_227; // @[FFT.scala 34:12]
  wire [31:0] _GEN_228; // @[FFT.scala 34:12]
  wire [31:0] _GEN_229; // @[FFT.scala 34:12]
  wire [31:0] _GEN_230; // @[FFT.scala 34:12]
  wire [31:0] _GEN_231; // @[FFT.scala 34:12]
  wire [31:0] _GEN_232; // @[FFT.scala 34:12]
  wire [31:0] _GEN_233; // @[FFT.scala 34:12]
  wire [31:0] _GEN_234; // @[FFT.scala 34:12]
  wire [31:0] _GEN_235; // @[FFT.scala 34:12]
  wire [31:0] _GEN_236; // @[FFT.scala 34:12]
  wire [31:0] _GEN_237; // @[FFT.scala 34:12]
  wire [31:0] _GEN_238; // @[FFT.scala 34:12]
  wire [31:0] _GEN_239; // @[FFT.scala 34:12]
  wire [31:0] _GEN_240; // @[FFT.scala 34:12]
  wire [31:0] _GEN_241; // @[FFT.scala 34:12]
  wire [31:0] _GEN_242; // @[FFT.scala 34:12]
  wire [31:0] _GEN_243; // @[FFT.scala 34:12]
  wire [31:0] _GEN_244; // @[FFT.scala 34:12]
  wire [31:0] _GEN_245; // @[FFT.scala 34:12]
  wire [31:0] _GEN_246; // @[FFT.scala 34:12]
  wire [31:0] _GEN_247; // @[FFT.scala 34:12]
  wire [31:0] _GEN_248; // @[FFT.scala 34:12]
  wire [31:0] _GEN_249; // @[FFT.scala 34:12]
  wire [31:0] _GEN_250; // @[FFT.scala 34:12]
  wire [31:0] _GEN_251; // @[FFT.scala 34:12]
  wire [31:0] _GEN_252; // @[FFT.scala 34:12]
  wire [31:0] _GEN_253; // @[FFT.scala 34:12]
  wire [31:0] _GEN_254; // @[FFT.scala 34:12]
  wire [31:0] _GEN_255; // @[FFT.scala 34:12]
  wire [31:0] _GEN_256; // @[FFT.scala 34:12]
  wire [31:0] _GEN_257; // @[FFT.scala 34:12]
  wire [31:0] _GEN_258; // @[FFT.scala 34:12]
  wire [31:0] _GEN_259; // @[FFT.scala 34:12]
  wire [31:0] _GEN_260; // @[FFT.scala 34:12]
  wire [31:0] _GEN_261; // @[FFT.scala 34:12]
  wire [31:0] _GEN_262; // @[FFT.scala 34:12]
  wire [31:0] _GEN_263; // @[FFT.scala 34:12]
  wire [31:0] _GEN_264; // @[FFT.scala 34:12]
  wire [31:0] _GEN_265; // @[FFT.scala 34:12]
  wire [31:0] _GEN_266; // @[FFT.scala 34:12]
  wire [31:0] _GEN_267; // @[FFT.scala 34:12]
  wire [31:0] _GEN_268; // @[FFT.scala 34:12]
  wire [31:0] _GEN_269; // @[FFT.scala 34:12]
  wire [31:0] _GEN_270; // @[FFT.scala 34:12]
  wire [31:0] _GEN_271; // @[FFT.scala 34:12]
  wire [31:0] _GEN_272; // @[FFT.scala 34:12]
  wire [31:0] _GEN_273; // @[FFT.scala 34:12]
  wire [31:0] _GEN_274; // @[FFT.scala 34:12]
  wire [31:0] _GEN_275; // @[FFT.scala 34:12]
  wire [31:0] _GEN_276; // @[FFT.scala 34:12]
  wire [31:0] _GEN_277; // @[FFT.scala 34:12]
  wire [31:0] _GEN_278; // @[FFT.scala 34:12]
  wire [31:0] _GEN_279; // @[FFT.scala 34:12]
  wire [31:0] _GEN_280; // @[FFT.scala 34:12]
  wire [31:0] _GEN_281; // @[FFT.scala 34:12]
  wire [31:0] _GEN_282; // @[FFT.scala 34:12]
  wire [31:0] _GEN_283; // @[FFT.scala 34:12]
  wire [31:0] _GEN_284; // @[FFT.scala 34:12]
  wire [31:0] _GEN_285; // @[FFT.scala 34:12]
  wire [31:0] _GEN_286; // @[FFT.scala 34:12]
  wire [31:0] _GEN_287; // @[FFT.scala 34:12]
  wire [31:0] _GEN_288; // @[FFT.scala 34:12]
  wire [31:0] _GEN_289; // @[FFT.scala 34:12]
  wire [31:0] _GEN_290; // @[FFT.scala 34:12]
  wire [31:0] _GEN_291; // @[FFT.scala 34:12]
  wire [31:0] _GEN_292; // @[FFT.scala 34:12]
  wire [31:0] _GEN_293; // @[FFT.scala 34:12]
  wire [31:0] _GEN_294; // @[FFT.scala 34:12]
  wire [31:0] _GEN_295; // @[FFT.scala 34:12]
  wire [31:0] _GEN_296; // @[FFT.scala 34:12]
  wire [31:0] _GEN_297; // @[FFT.scala 34:12]
  wire [31:0] _GEN_298; // @[FFT.scala 34:12]
  wire [31:0] _GEN_299; // @[FFT.scala 34:12]
  wire [31:0] _GEN_300; // @[FFT.scala 34:12]
  wire [31:0] _GEN_301; // @[FFT.scala 34:12]
  wire [31:0] _GEN_302; // @[FFT.scala 34:12]
  wire [31:0] _GEN_303; // @[FFT.scala 34:12]
  wire [31:0] _GEN_304; // @[FFT.scala 34:12]
  wire [31:0] _GEN_305; // @[FFT.scala 34:12]
  wire [31:0] _GEN_306; // @[FFT.scala 34:12]
  wire [31:0] _GEN_307; // @[FFT.scala 34:12]
  wire [31:0] _GEN_308; // @[FFT.scala 34:12]
  wire [31:0] _GEN_309; // @[FFT.scala 34:12]
  wire [31:0] _GEN_310; // @[FFT.scala 34:12]
  wire [31:0] _GEN_311; // @[FFT.scala 34:12]
  wire [31:0] _GEN_312; // @[FFT.scala 34:12]
  wire [31:0] _GEN_313; // @[FFT.scala 34:12]
  wire [31:0] _GEN_314; // @[FFT.scala 34:12]
  wire [31:0] _GEN_315; // @[FFT.scala 34:12]
  wire [31:0] _GEN_316; // @[FFT.scala 34:12]
  wire [31:0] _GEN_317; // @[FFT.scala 34:12]
  wire [31:0] _GEN_318; // @[FFT.scala 34:12]
  wire [31:0] _GEN_319; // @[FFT.scala 34:12]
  wire [31:0] _GEN_320; // @[FFT.scala 34:12]
  wire [31:0] _GEN_321; // @[FFT.scala 34:12]
  wire [31:0] _GEN_322; // @[FFT.scala 34:12]
  wire [31:0] _GEN_323; // @[FFT.scala 34:12]
  wire [31:0] _GEN_324; // @[FFT.scala 34:12]
  wire [31:0] _GEN_325; // @[FFT.scala 34:12]
  wire [31:0] _GEN_326; // @[FFT.scala 34:12]
  wire [31:0] _GEN_327; // @[FFT.scala 34:12]
  wire [31:0] _GEN_328; // @[FFT.scala 34:12]
  wire [31:0] _GEN_329; // @[FFT.scala 34:12]
  wire [31:0] _GEN_330; // @[FFT.scala 34:12]
  wire [31:0] _GEN_331; // @[FFT.scala 34:12]
  wire [31:0] _GEN_332; // @[FFT.scala 34:12]
  wire [31:0] _GEN_333; // @[FFT.scala 34:12]
  wire [31:0] _GEN_334; // @[FFT.scala 34:12]
  wire [31:0] _GEN_335; // @[FFT.scala 34:12]
  wire [31:0] _GEN_336; // @[FFT.scala 34:12]
  wire [31:0] _GEN_337; // @[FFT.scala 34:12]
  wire [31:0] _GEN_338; // @[FFT.scala 34:12]
  wire [31:0] _GEN_339; // @[FFT.scala 34:12]
  wire [31:0] _GEN_340; // @[FFT.scala 34:12]
  wire [31:0] _GEN_341; // @[FFT.scala 34:12]
  wire [31:0] _GEN_342; // @[FFT.scala 34:12]
  wire [31:0] _GEN_343; // @[FFT.scala 34:12]
  wire [31:0] _GEN_344; // @[FFT.scala 34:12]
  wire [31:0] _GEN_345; // @[FFT.scala 34:12]
  wire [31:0] _GEN_346; // @[FFT.scala 34:12]
  wire [31:0] _GEN_347; // @[FFT.scala 34:12]
  wire [31:0] _GEN_348; // @[FFT.scala 34:12]
  wire [31:0] _GEN_349; // @[FFT.scala 34:12]
  wire [31:0] _GEN_350; // @[FFT.scala 34:12]
  wire [31:0] _GEN_351; // @[FFT.scala 34:12]
  wire [31:0] _GEN_352; // @[FFT.scala 34:12]
  wire [31:0] _GEN_353; // @[FFT.scala 34:12]
  wire [31:0] _GEN_354; // @[FFT.scala 34:12]
  wire [31:0] _GEN_355; // @[FFT.scala 34:12]
  wire [31:0] _GEN_356; // @[FFT.scala 34:12]
  wire [31:0] _GEN_357; // @[FFT.scala 34:12]
  wire [31:0] _GEN_358; // @[FFT.scala 34:12]
  wire [31:0] _GEN_359; // @[FFT.scala 34:12]
  wire [31:0] _GEN_360; // @[FFT.scala 34:12]
  wire [31:0] _GEN_361; // @[FFT.scala 34:12]
  wire [31:0] _GEN_362; // @[FFT.scala 34:12]
  wire [31:0] _GEN_363; // @[FFT.scala 34:12]
  wire [31:0] _GEN_364; // @[FFT.scala 34:12]
  wire [31:0] _GEN_365; // @[FFT.scala 34:12]
  wire [31:0] _GEN_366; // @[FFT.scala 34:12]
  wire [31:0] _GEN_367; // @[FFT.scala 34:12]
  wire [31:0] _GEN_368; // @[FFT.scala 34:12]
  wire [31:0] _GEN_369; // @[FFT.scala 34:12]
  wire [31:0] _GEN_370; // @[FFT.scala 34:12]
  wire [31:0] _GEN_371; // @[FFT.scala 34:12]
  wire [31:0] _GEN_372; // @[FFT.scala 34:12]
  wire [31:0] _GEN_373; // @[FFT.scala 34:12]
  wire [31:0] _GEN_374; // @[FFT.scala 34:12]
  wire [31:0] _GEN_375; // @[FFT.scala 34:12]
  wire [31:0] _GEN_376; // @[FFT.scala 34:12]
  wire [31:0] _GEN_377; // @[FFT.scala 34:12]
  wire [31:0] _GEN_378; // @[FFT.scala 34:12]
  wire [31:0] _GEN_379; // @[FFT.scala 34:12]
  wire [31:0] _GEN_380; // @[FFT.scala 34:12]
  wire [31:0] _GEN_381; // @[FFT.scala 34:12]
  wire [31:0] _GEN_382; // @[FFT.scala 34:12]
  wire [31:0] _GEN_383; // @[FFT.scala 34:12]
  wire [31:0] _GEN_384; // @[FFT.scala 34:12]
  wire [31:0] _GEN_385; // @[FFT.scala 34:12]
  wire [31:0] _GEN_386; // @[FFT.scala 34:12]
  wire [31:0] _GEN_387; // @[FFT.scala 34:12]
  wire [31:0] _GEN_388; // @[FFT.scala 34:12]
  wire [31:0] _GEN_389; // @[FFT.scala 34:12]
  wire [31:0] _GEN_390; // @[FFT.scala 34:12]
  wire [31:0] _GEN_391; // @[FFT.scala 34:12]
  wire [31:0] _GEN_392; // @[FFT.scala 34:12]
  wire [31:0] _GEN_393; // @[FFT.scala 34:12]
  wire [31:0] _GEN_394; // @[FFT.scala 34:12]
  wire [31:0] _GEN_395; // @[FFT.scala 34:12]
  wire [31:0] _GEN_396; // @[FFT.scala 34:12]
  wire [31:0] _GEN_397; // @[FFT.scala 34:12]
  wire [31:0] _GEN_398; // @[FFT.scala 34:12]
  wire [31:0] _GEN_399; // @[FFT.scala 34:12]
  wire [31:0] _GEN_400; // @[FFT.scala 34:12]
  wire [31:0] _GEN_401; // @[FFT.scala 34:12]
  wire [31:0] _GEN_402; // @[FFT.scala 34:12]
  wire [31:0] _GEN_403; // @[FFT.scala 34:12]
  wire [31:0] _GEN_404; // @[FFT.scala 34:12]
  wire [31:0] _GEN_405; // @[FFT.scala 34:12]
  wire [31:0] _GEN_406; // @[FFT.scala 34:12]
  wire [31:0] _GEN_407; // @[FFT.scala 34:12]
  wire [31:0] _GEN_408; // @[FFT.scala 34:12]
  wire [31:0] _GEN_409; // @[FFT.scala 34:12]
  wire [31:0] _GEN_410; // @[FFT.scala 34:12]
  wire [31:0] _GEN_411; // @[FFT.scala 34:12]
  wire [31:0] _GEN_412; // @[FFT.scala 34:12]
  wire [31:0] _GEN_413; // @[FFT.scala 34:12]
  wire [31:0] _GEN_414; // @[FFT.scala 34:12]
  wire [31:0] _GEN_415; // @[FFT.scala 34:12]
  wire [31:0] _GEN_416; // @[FFT.scala 34:12]
  wire [31:0] _GEN_417; // @[FFT.scala 34:12]
  wire [31:0] _GEN_418; // @[FFT.scala 34:12]
  wire [31:0] _GEN_419; // @[FFT.scala 34:12]
  wire [31:0] _GEN_420; // @[FFT.scala 34:12]
  wire [31:0] _GEN_421; // @[FFT.scala 34:12]
  wire [31:0] _GEN_422; // @[FFT.scala 34:12]
  wire [31:0] _GEN_423; // @[FFT.scala 34:12]
  wire [31:0] _GEN_424; // @[FFT.scala 34:12]
  wire [31:0] _GEN_425; // @[FFT.scala 34:12]
  wire [31:0] _GEN_426; // @[FFT.scala 34:12]
  wire [31:0] _GEN_427; // @[FFT.scala 34:12]
  wire [31:0] _GEN_428; // @[FFT.scala 34:12]
  wire [31:0] _GEN_429; // @[FFT.scala 34:12]
  wire [31:0] _GEN_430; // @[FFT.scala 34:12]
  wire [31:0] _GEN_431; // @[FFT.scala 34:12]
  wire [31:0] _GEN_432; // @[FFT.scala 34:12]
  wire [31:0] _GEN_433; // @[FFT.scala 34:12]
  wire [31:0] _GEN_434; // @[FFT.scala 34:12]
  wire [31:0] _GEN_435; // @[FFT.scala 34:12]
  wire [31:0] _GEN_436; // @[FFT.scala 34:12]
  wire [31:0] _GEN_437; // @[FFT.scala 34:12]
  wire [31:0] _GEN_438; // @[FFT.scala 34:12]
  wire [31:0] _GEN_439; // @[FFT.scala 34:12]
  wire [31:0] _GEN_440; // @[FFT.scala 34:12]
  wire [31:0] _GEN_441; // @[FFT.scala 34:12]
  wire [31:0] _GEN_442; // @[FFT.scala 34:12]
  wire [31:0] _GEN_443; // @[FFT.scala 34:12]
  wire [31:0] _GEN_444; // @[FFT.scala 34:12]
  wire [31:0] _GEN_445; // @[FFT.scala 34:12]
  wire [31:0] _GEN_446; // @[FFT.scala 34:12]
  wire [31:0] _GEN_447; // @[FFT.scala 34:12]
  wire [31:0] _GEN_448; // @[FFT.scala 34:12]
  wire [31:0] _GEN_449; // @[FFT.scala 34:12]
  wire [31:0] _GEN_450; // @[FFT.scala 34:12]
  wire [31:0] _GEN_451; // @[FFT.scala 34:12]
  wire [31:0] _GEN_452; // @[FFT.scala 34:12]
  wire [31:0] _GEN_453; // @[FFT.scala 34:12]
  wire [31:0] _GEN_454; // @[FFT.scala 34:12]
  wire [31:0] _GEN_455; // @[FFT.scala 34:12]
  wire [31:0] _GEN_456; // @[FFT.scala 34:12]
  wire [31:0] _GEN_457; // @[FFT.scala 34:12]
  wire [31:0] _GEN_458; // @[FFT.scala 34:12]
  wire [31:0] _GEN_459; // @[FFT.scala 34:12]
  wire [31:0] _GEN_460; // @[FFT.scala 34:12]
  wire [31:0] _GEN_461; // @[FFT.scala 34:12]
  wire [31:0] _GEN_462; // @[FFT.scala 34:12]
  wire [31:0] _GEN_463; // @[FFT.scala 34:12]
  wire [31:0] _GEN_464; // @[FFT.scala 34:12]
  wire [31:0] _GEN_465; // @[FFT.scala 34:12]
  wire [31:0] _GEN_466; // @[FFT.scala 34:12]
  wire [31:0] _GEN_467; // @[FFT.scala 34:12]
  wire [31:0] _GEN_468; // @[FFT.scala 34:12]
  wire [31:0] _GEN_469; // @[FFT.scala 34:12]
  wire [31:0] _GEN_470; // @[FFT.scala 34:12]
  wire [31:0] _GEN_471; // @[FFT.scala 34:12]
  wire [31:0] _GEN_472; // @[FFT.scala 34:12]
  wire [31:0] _GEN_473; // @[FFT.scala 34:12]
  wire [31:0] _GEN_474; // @[FFT.scala 34:12]
  wire [31:0] _GEN_475; // @[FFT.scala 34:12]
  wire [31:0] _GEN_476; // @[FFT.scala 34:12]
  wire [31:0] _GEN_477; // @[FFT.scala 34:12]
  wire [31:0] _GEN_478; // @[FFT.scala 34:12]
  wire [31:0] _GEN_479; // @[FFT.scala 34:12]
  wire [31:0] _GEN_480; // @[FFT.scala 34:12]
  wire [31:0] _GEN_481; // @[FFT.scala 34:12]
  wire [31:0] _GEN_482; // @[FFT.scala 34:12]
  wire [31:0] _GEN_483; // @[FFT.scala 34:12]
  wire [31:0] _GEN_484; // @[FFT.scala 34:12]
  wire [31:0] _GEN_485; // @[FFT.scala 34:12]
  wire [31:0] _GEN_486; // @[FFT.scala 34:12]
  wire [31:0] _GEN_487; // @[FFT.scala 34:12]
  wire [31:0] _GEN_488; // @[FFT.scala 34:12]
  wire [31:0] _GEN_489; // @[FFT.scala 34:12]
  wire [31:0] _GEN_490; // @[FFT.scala 34:12]
  wire [31:0] _GEN_491; // @[FFT.scala 34:12]
  wire [31:0] _GEN_492; // @[FFT.scala 34:12]
  wire [31:0] _GEN_493; // @[FFT.scala 34:12]
  wire [31:0] _GEN_494; // @[FFT.scala 34:12]
  wire [31:0] _GEN_495; // @[FFT.scala 34:12]
  wire [31:0] _GEN_496; // @[FFT.scala 34:12]
  wire [31:0] _GEN_497; // @[FFT.scala 34:12]
  wire [31:0] _GEN_498; // @[FFT.scala 34:12]
  wire [31:0] _GEN_499; // @[FFT.scala 34:12]
  wire [31:0] _GEN_500; // @[FFT.scala 34:12]
  wire [31:0] _GEN_501; // @[FFT.scala 34:12]
  wire [31:0] _GEN_502; // @[FFT.scala 34:12]
  wire [31:0] _GEN_503; // @[FFT.scala 34:12]
  wire [31:0] _GEN_504; // @[FFT.scala 34:12]
  wire [31:0] _GEN_505; // @[FFT.scala 34:12]
  wire [31:0] _GEN_506; // @[FFT.scala 34:12]
  wire [31:0] _GEN_507; // @[FFT.scala 34:12]
  wire [31:0] _GEN_508; // @[FFT.scala 34:12]
  wire [31:0] _GEN_509; // @[FFT.scala 34:12]
  wire [31:0] _GEN_510; // @[FFT.scala 34:12]
  wire [31:0] _GEN_511; // @[FFT.scala 34:12]
  wire [31:0] _GEN_514; // @[FFT.scala 35:12]
  wire [31:0] _GEN_515; // @[FFT.scala 35:12]
  wire [31:0] _GEN_516; // @[FFT.scala 35:12]
  wire [31:0] _GEN_517; // @[FFT.scala 35:12]
  wire [31:0] _GEN_518; // @[FFT.scala 35:12]
  wire [31:0] _GEN_519; // @[FFT.scala 35:12]
  wire [31:0] _GEN_520; // @[FFT.scala 35:12]
  wire [31:0] _GEN_521; // @[FFT.scala 35:12]
  wire [31:0] _GEN_522; // @[FFT.scala 35:12]
  wire [31:0] _GEN_523; // @[FFT.scala 35:12]
  wire [31:0] _GEN_524; // @[FFT.scala 35:12]
  wire [31:0] _GEN_525; // @[FFT.scala 35:12]
  wire [31:0] _GEN_526; // @[FFT.scala 35:12]
  wire [31:0] _GEN_527; // @[FFT.scala 35:12]
  wire [31:0] _GEN_528; // @[FFT.scala 35:12]
  wire [31:0] _GEN_529; // @[FFT.scala 35:12]
  wire [31:0] _GEN_530; // @[FFT.scala 35:12]
  wire [31:0] _GEN_531; // @[FFT.scala 35:12]
  wire [31:0] _GEN_532; // @[FFT.scala 35:12]
  wire [31:0] _GEN_533; // @[FFT.scala 35:12]
  wire [31:0] _GEN_534; // @[FFT.scala 35:12]
  wire [31:0] _GEN_535; // @[FFT.scala 35:12]
  wire [31:0] _GEN_536; // @[FFT.scala 35:12]
  wire [31:0] _GEN_537; // @[FFT.scala 35:12]
  wire [31:0] _GEN_538; // @[FFT.scala 35:12]
  wire [31:0] _GEN_539; // @[FFT.scala 35:12]
  wire [31:0] _GEN_540; // @[FFT.scala 35:12]
  wire [31:0] _GEN_541; // @[FFT.scala 35:12]
  wire [31:0] _GEN_542; // @[FFT.scala 35:12]
  wire [31:0] _GEN_543; // @[FFT.scala 35:12]
  wire [31:0] _GEN_544; // @[FFT.scala 35:12]
  wire [31:0] _GEN_545; // @[FFT.scala 35:12]
  wire [31:0] _GEN_546; // @[FFT.scala 35:12]
  wire [31:0] _GEN_547; // @[FFT.scala 35:12]
  wire [31:0] _GEN_548; // @[FFT.scala 35:12]
  wire [31:0] _GEN_549; // @[FFT.scala 35:12]
  wire [31:0] _GEN_550; // @[FFT.scala 35:12]
  wire [31:0] _GEN_551; // @[FFT.scala 35:12]
  wire [31:0] _GEN_552; // @[FFT.scala 35:12]
  wire [31:0] _GEN_553; // @[FFT.scala 35:12]
  wire [31:0] _GEN_554; // @[FFT.scala 35:12]
  wire [31:0] _GEN_555; // @[FFT.scala 35:12]
  wire [31:0] _GEN_556; // @[FFT.scala 35:12]
  wire [31:0] _GEN_557; // @[FFT.scala 35:12]
  wire [31:0] _GEN_558; // @[FFT.scala 35:12]
  wire [31:0] _GEN_559; // @[FFT.scala 35:12]
  wire [31:0] _GEN_560; // @[FFT.scala 35:12]
  wire [31:0] _GEN_561; // @[FFT.scala 35:12]
  wire [31:0] _GEN_562; // @[FFT.scala 35:12]
  wire [31:0] _GEN_563; // @[FFT.scala 35:12]
  wire [31:0] _GEN_564; // @[FFT.scala 35:12]
  wire [31:0] _GEN_565; // @[FFT.scala 35:12]
  wire [31:0] _GEN_566; // @[FFT.scala 35:12]
  wire [31:0] _GEN_567; // @[FFT.scala 35:12]
  wire [31:0] _GEN_568; // @[FFT.scala 35:12]
  wire [31:0] _GEN_569; // @[FFT.scala 35:12]
  wire [31:0] _GEN_570; // @[FFT.scala 35:12]
  wire [31:0] _GEN_571; // @[FFT.scala 35:12]
  wire [31:0] _GEN_572; // @[FFT.scala 35:12]
  wire [31:0] _GEN_573; // @[FFT.scala 35:12]
  wire [31:0] _GEN_574; // @[FFT.scala 35:12]
  wire [31:0] _GEN_575; // @[FFT.scala 35:12]
  wire [31:0] _GEN_576; // @[FFT.scala 35:12]
  wire [31:0] _GEN_577; // @[FFT.scala 35:12]
  wire [31:0] _GEN_578; // @[FFT.scala 35:12]
  wire [31:0] _GEN_579; // @[FFT.scala 35:12]
  wire [31:0] _GEN_580; // @[FFT.scala 35:12]
  wire [31:0] _GEN_581; // @[FFT.scala 35:12]
  wire [31:0] _GEN_582; // @[FFT.scala 35:12]
  wire [31:0] _GEN_583; // @[FFT.scala 35:12]
  wire [31:0] _GEN_584; // @[FFT.scala 35:12]
  wire [31:0] _GEN_585; // @[FFT.scala 35:12]
  wire [31:0] _GEN_586; // @[FFT.scala 35:12]
  wire [31:0] _GEN_587; // @[FFT.scala 35:12]
  wire [31:0] _GEN_588; // @[FFT.scala 35:12]
  wire [31:0] _GEN_589; // @[FFT.scala 35:12]
  wire [31:0] _GEN_590; // @[FFT.scala 35:12]
  wire [31:0] _GEN_591; // @[FFT.scala 35:12]
  wire [31:0] _GEN_592; // @[FFT.scala 35:12]
  wire [31:0] _GEN_593; // @[FFT.scala 35:12]
  wire [31:0] _GEN_594; // @[FFT.scala 35:12]
  wire [31:0] _GEN_595; // @[FFT.scala 35:12]
  wire [31:0] _GEN_596; // @[FFT.scala 35:12]
  wire [31:0] _GEN_597; // @[FFT.scala 35:12]
  wire [31:0] _GEN_598; // @[FFT.scala 35:12]
  wire [31:0] _GEN_599; // @[FFT.scala 35:12]
  wire [31:0] _GEN_600; // @[FFT.scala 35:12]
  wire [31:0] _GEN_601; // @[FFT.scala 35:12]
  wire [31:0] _GEN_602; // @[FFT.scala 35:12]
  wire [31:0] _GEN_603; // @[FFT.scala 35:12]
  wire [31:0] _GEN_604; // @[FFT.scala 35:12]
  wire [31:0] _GEN_605; // @[FFT.scala 35:12]
  wire [31:0] _GEN_606; // @[FFT.scala 35:12]
  wire [31:0] _GEN_607; // @[FFT.scala 35:12]
  wire [31:0] _GEN_608; // @[FFT.scala 35:12]
  wire [31:0] _GEN_609; // @[FFT.scala 35:12]
  wire [31:0] _GEN_610; // @[FFT.scala 35:12]
  wire [31:0] _GEN_611; // @[FFT.scala 35:12]
  wire [31:0] _GEN_612; // @[FFT.scala 35:12]
  wire [31:0] _GEN_613; // @[FFT.scala 35:12]
  wire [31:0] _GEN_614; // @[FFT.scala 35:12]
  wire [31:0] _GEN_615; // @[FFT.scala 35:12]
  wire [31:0] _GEN_616; // @[FFT.scala 35:12]
  wire [31:0] _GEN_617; // @[FFT.scala 35:12]
  wire [31:0] _GEN_618; // @[FFT.scala 35:12]
  wire [31:0] _GEN_619; // @[FFT.scala 35:12]
  wire [31:0] _GEN_620; // @[FFT.scala 35:12]
  wire [31:0] _GEN_621; // @[FFT.scala 35:12]
  wire [31:0] _GEN_622; // @[FFT.scala 35:12]
  wire [31:0] _GEN_623; // @[FFT.scala 35:12]
  wire [31:0] _GEN_624; // @[FFT.scala 35:12]
  wire [31:0] _GEN_625; // @[FFT.scala 35:12]
  wire [31:0] _GEN_626; // @[FFT.scala 35:12]
  wire [31:0] _GEN_627; // @[FFT.scala 35:12]
  wire [31:0] _GEN_628; // @[FFT.scala 35:12]
  wire [31:0] _GEN_629; // @[FFT.scala 35:12]
  wire [31:0] _GEN_630; // @[FFT.scala 35:12]
  wire [31:0] _GEN_631; // @[FFT.scala 35:12]
  wire [31:0] _GEN_632; // @[FFT.scala 35:12]
  wire [31:0] _GEN_633; // @[FFT.scala 35:12]
  wire [31:0] _GEN_634; // @[FFT.scala 35:12]
  wire [31:0] _GEN_635; // @[FFT.scala 35:12]
  wire [31:0] _GEN_636; // @[FFT.scala 35:12]
  wire [31:0] _GEN_637; // @[FFT.scala 35:12]
  wire [31:0] _GEN_638; // @[FFT.scala 35:12]
  wire [31:0] _GEN_639; // @[FFT.scala 35:12]
  wire [31:0] _GEN_640; // @[FFT.scala 35:12]
  wire [31:0] _GEN_641; // @[FFT.scala 35:12]
  wire [31:0] _GEN_642; // @[FFT.scala 35:12]
  wire [31:0] _GEN_643; // @[FFT.scala 35:12]
  wire [31:0] _GEN_644; // @[FFT.scala 35:12]
  wire [31:0] _GEN_645; // @[FFT.scala 35:12]
  wire [31:0] _GEN_646; // @[FFT.scala 35:12]
  wire [31:0] _GEN_647; // @[FFT.scala 35:12]
  wire [31:0] _GEN_648; // @[FFT.scala 35:12]
  wire [31:0] _GEN_649; // @[FFT.scala 35:12]
  wire [31:0] _GEN_650; // @[FFT.scala 35:12]
  wire [31:0] _GEN_651; // @[FFT.scala 35:12]
  wire [31:0] _GEN_652; // @[FFT.scala 35:12]
  wire [31:0] _GEN_653; // @[FFT.scala 35:12]
  wire [31:0] _GEN_654; // @[FFT.scala 35:12]
  wire [31:0] _GEN_655; // @[FFT.scala 35:12]
  wire [31:0] _GEN_656; // @[FFT.scala 35:12]
  wire [31:0] _GEN_657; // @[FFT.scala 35:12]
  wire [31:0] _GEN_658; // @[FFT.scala 35:12]
  wire [31:0] _GEN_659; // @[FFT.scala 35:12]
  wire [31:0] _GEN_660; // @[FFT.scala 35:12]
  wire [31:0] _GEN_661; // @[FFT.scala 35:12]
  wire [31:0] _GEN_662; // @[FFT.scala 35:12]
  wire [31:0] _GEN_663; // @[FFT.scala 35:12]
  wire [31:0] _GEN_664; // @[FFT.scala 35:12]
  wire [31:0] _GEN_665; // @[FFT.scala 35:12]
  wire [31:0] _GEN_666; // @[FFT.scala 35:12]
  wire [31:0] _GEN_667; // @[FFT.scala 35:12]
  wire [31:0] _GEN_668; // @[FFT.scala 35:12]
  wire [31:0] _GEN_669; // @[FFT.scala 35:12]
  wire [31:0] _GEN_670; // @[FFT.scala 35:12]
  wire [31:0] _GEN_671; // @[FFT.scala 35:12]
  wire [31:0] _GEN_672; // @[FFT.scala 35:12]
  wire [31:0] _GEN_673; // @[FFT.scala 35:12]
  wire [31:0] _GEN_674; // @[FFT.scala 35:12]
  wire [31:0] _GEN_675; // @[FFT.scala 35:12]
  wire [31:0] _GEN_676; // @[FFT.scala 35:12]
  wire [31:0] _GEN_677; // @[FFT.scala 35:12]
  wire [31:0] _GEN_678; // @[FFT.scala 35:12]
  wire [31:0] _GEN_679; // @[FFT.scala 35:12]
  wire [31:0] _GEN_680; // @[FFT.scala 35:12]
  wire [31:0] _GEN_681; // @[FFT.scala 35:12]
  wire [31:0] _GEN_682; // @[FFT.scala 35:12]
  wire [31:0] _GEN_683; // @[FFT.scala 35:12]
  wire [31:0] _GEN_684; // @[FFT.scala 35:12]
  wire [31:0] _GEN_685; // @[FFT.scala 35:12]
  wire [31:0] _GEN_686; // @[FFT.scala 35:12]
  wire [31:0] _GEN_687; // @[FFT.scala 35:12]
  wire [31:0] _GEN_688; // @[FFT.scala 35:12]
  wire [31:0] _GEN_689; // @[FFT.scala 35:12]
  wire [31:0] _GEN_690; // @[FFT.scala 35:12]
  wire [31:0] _GEN_691; // @[FFT.scala 35:12]
  wire [31:0] _GEN_692; // @[FFT.scala 35:12]
  wire [31:0] _GEN_693; // @[FFT.scala 35:12]
  wire [31:0] _GEN_694; // @[FFT.scala 35:12]
  wire [31:0] _GEN_695; // @[FFT.scala 35:12]
  wire [31:0] _GEN_696; // @[FFT.scala 35:12]
  wire [31:0] _GEN_697; // @[FFT.scala 35:12]
  wire [31:0] _GEN_698; // @[FFT.scala 35:12]
  wire [31:0] _GEN_699; // @[FFT.scala 35:12]
  wire [31:0] _GEN_700; // @[FFT.scala 35:12]
  wire [31:0] _GEN_701; // @[FFT.scala 35:12]
  wire [31:0] _GEN_702; // @[FFT.scala 35:12]
  wire [31:0] _GEN_703; // @[FFT.scala 35:12]
  wire [31:0] _GEN_704; // @[FFT.scala 35:12]
  wire [31:0] _GEN_705; // @[FFT.scala 35:12]
  wire [31:0] _GEN_706; // @[FFT.scala 35:12]
  wire [31:0] _GEN_707; // @[FFT.scala 35:12]
  wire [31:0] _GEN_708; // @[FFT.scala 35:12]
  wire [31:0] _GEN_709; // @[FFT.scala 35:12]
  wire [31:0] _GEN_710; // @[FFT.scala 35:12]
  wire [31:0] _GEN_711; // @[FFT.scala 35:12]
  wire [31:0] _GEN_712; // @[FFT.scala 35:12]
  wire [31:0] _GEN_713; // @[FFT.scala 35:12]
  wire [31:0] _GEN_714; // @[FFT.scala 35:12]
  wire [31:0] _GEN_715; // @[FFT.scala 35:12]
  wire [31:0] _GEN_716; // @[FFT.scala 35:12]
  wire [31:0] _GEN_717; // @[FFT.scala 35:12]
  wire [31:0] _GEN_718; // @[FFT.scala 35:12]
  wire [31:0] _GEN_719; // @[FFT.scala 35:12]
  wire [31:0] _GEN_720; // @[FFT.scala 35:12]
  wire [31:0] _GEN_721; // @[FFT.scala 35:12]
  wire [31:0] _GEN_722; // @[FFT.scala 35:12]
  wire [31:0] _GEN_723; // @[FFT.scala 35:12]
  wire [31:0] _GEN_724; // @[FFT.scala 35:12]
  wire [31:0] _GEN_725; // @[FFT.scala 35:12]
  wire [31:0] _GEN_726; // @[FFT.scala 35:12]
  wire [31:0] _GEN_727; // @[FFT.scala 35:12]
  wire [31:0] _GEN_728; // @[FFT.scala 35:12]
  wire [31:0] _GEN_729; // @[FFT.scala 35:12]
  wire [31:0] _GEN_730; // @[FFT.scala 35:12]
  wire [31:0] _GEN_731; // @[FFT.scala 35:12]
  wire [31:0] _GEN_732; // @[FFT.scala 35:12]
  wire [31:0] _GEN_733; // @[FFT.scala 35:12]
  wire [31:0] _GEN_734; // @[FFT.scala 35:12]
  wire [31:0] _GEN_735; // @[FFT.scala 35:12]
  wire [31:0] _GEN_736; // @[FFT.scala 35:12]
  wire [31:0] _GEN_737; // @[FFT.scala 35:12]
  wire [31:0] _GEN_738; // @[FFT.scala 35:12]
  wire [31:0] _GEN_739; // @[FFT.scala 35:12]
  wire [31:0] _GEN_740; // @[FFT.scala 35:12]
  wire [31:0] _GEN_741; // @[FFT.scala 35:12]
  wire [31:0] _GEN_742; // @[FFT.scala 35:12]
  wire [31:0] _GEN_743; // @[FFT.scala 35:12]
  wire [31:0] _GEN_744; // @[FFT.scala 35:12]
  wire [31:0] _GEN_745; // @[FFT.scala 35:12]
  wire [31:0] _GEN_746; // @[FFT.scala 35:12]
  wire [31:0] _GEN_747; // @[FFT.scala 35:12]
  wire [31:0] _GEN_748; // @[FFT.scala 35:12]
  wire [31:0] _GEN_749; // @[FFT.scala 35:12]
  wire [31:0] _GEN_750; // @[FFT.scala 35:12]
  wire [31:0] _GEN_751; // @[FFT.scala 35:12]
  wire [31:0] _GEN_752; // @[FFT.scala 35:12]
  wire [31:0] _GEN_753; // @[FFT.scala 35:12]
  wire [31:0] _GEN_754; // @[FFT.scala 35:12]
  wire [31:0] _GEN_755; // @[FFT.scala 35:12]
  wire [31:0] _GEN_756; // @[FFT.scala 35:12]
  wire [31:0] _GEN_757; // @[FFT.scala 35:12]
  wire [31:0] _GEN_758; // @[FFT.scala 35:12]
  wire [31:0] _GEN_759; // @[FFT.scala 35:12]
  wire [31:0] _GEN_760; // @[FFT.scala 35:12]
  wire [31:0] _GEN_761; // @[FFT.scala 35:12]
  wire [31:0] _GEN_762; // @[FFT.scala 35:12]
  wire [31:0] _GEN_763; // @[FFT.scala 35:12]
  wire [31:0] _GEN_764; // @[FFT.scala 35:12]
  wire [31:0] _GEN_765; // @[FFT.scala 35:12]
  wire [31:0] _GEN_766; // @[FFT.scala 35:12]
  wire [31:0] _GEN_767; // @[FFT.scala 35:12]
  wire [31:0] _GEN_768; // @[FFT.scala 35:12]
  wire [31:0] _GEN_769; // @[FFT.scala 35:12]
  wire [31:0] _GEN_770; // @[FFT.scala 35:12]
  wire [31:0] _GEN_771; // @[FFT.scala 35:12]
  wire [31:0] _GEN_772; // @[FFT.scala 35:12]
  wire [31:0] _GEN_773; // @[FFT.scala 35:12]
  wire [31:0] _GEN_774; // @[FFT.scala 35:12]
  wire [31:0] _GEN_775; // @[FFT.scala 35:12]
  wire [31:0] _GEN_776; // @[FFT.scala 35:12]
  wire [31:0] _GEN_777; // @[FFT.scala 35:12]
  wire [31:0] _GEN_778; // @[FFT.scala 35:12]
  wire [31:0] _GEN_779; // @[FFT.scala 35:12]
  wire [31:0] _GEN_780; // @[FFT.scala 35:12]
  wire [31:0] _GEN_781; // @[FFT.scala 35:12]
  wire [31:0] _GEN_782; // @[FFT.scala 35:12]
  wire [31:0] _GEN_783; // @[FFT.scala 35:12]
  wire [31:0] _GEN_784; // @[FFT.scala 35:12]
  wire [31:0] _GEN_785; // @[FFT.scala 35:12]
  wire [31:0] _GEN_786; // @[FFT.scala 35:12]
  wire [31:0] _GEN_787; // @[FFT.scala 35:12]
  wire [31:0] _GEN_788; // @[FFT.scala 35:12]
  wire [31:0] _GEN_789; // @[FFT.scala 35:12]
  wire [31:0] _GEN_790; // @[FFT.scala 35:12]
  wire [31:0] _GEN_791; // @[FFT.scala 35:12]
  wire [31:0] _GEN_792; // @[FFT.scala 35:12]
  wire [31:0] _GEN_793; // @[FFT.scala 35:12]
  wire [31:0] _GEN_794; // @[FFT.scala 35:12]
  wire [31:0] _GEN_795; // @[FFT.scala 35:12]
  wire [31:0] _GEN_796; // @[FFT.scala 35:12]
  wire [31:0] _GEN_797; // @[FFT.scala 35:12]
  wire [31:0] _GEN_798; // @[FFT.scala 35:12]
  wire [31:0] _GEN_799; // @[FFT.scala 35:12]
  wire [31:0] _GEN_800; // @[FFT.scala 35:12]
  wire [31:0] _GEN_801; // @[FFT.scala 35:12]
  wire [31:0] _GEN_802; // @[FFT.scala 35:12]
  wire [31:0] _GEN_803; // @[FFT.scala 35:12]
  wire [31:0] _GEN_804; // @[FFT.scala 35:12]
  wire [31:0] _GEN_805; // @[FFT.scala 35:12]
  wire [31:0] _GEN_806; // @[FFT.scala 35:12]
  wire [31:0] _GEN_807; // @[FFT.scala 35:12]
  wire [31:0] _GEN_808; // @[FFT.scala 35:12]
  wire [31:0] _GEN_809; // @[FFT.scala 35:12]
  wire [31:0] _GEN_810; // @[FFT.scala 35:12]
  wire [31:0] _GEN_811; // @[FFT.scala 35:12]
  wire [31:0] _GEN_812; // @[FFT.scala 35:12]
  wire [31:0] _GEN_813; // @[FFT.scala 35:12]
  wire [31:0] _GEN_814; // @[FFT.scala 35:12]
  wire [31:0] _GEN_815; // @[FFT.scala 35:12]
  wire [31:0] _GEN_816; // @[FFT.scala 35:12]
  wire [31:0] _GEN_817; // @[FFT.scala 35:12]
  wire [31:0] _GEN_818; // @[FFT.scala 35:12]
  wire [31:0] _GEN_819; // @[FFT.scala 35:12]
  wire [31:0] _GEN_820; // @[FFT.scala 35:12]
  wire [31:0] _GEN_821; // @[FFT.scala 35:12]
  wire [31:0] _GEN_822; // @[FFT.scala 35:12]
  wire [31:0] _GEN_823; // @[FFT.scala 35:12]
  wire [31:0] _GEN_824; // @[FFT.scala 35:12]
  wire [31:0] _GEN_825; // @[FFT.scala 35:12]
  wire [31:0] _GEN_826; // @[FFT.scala 35:12]
  wire [31:0] _GEN_827; // @[FFT.scala 35:12]
  wire [31:0] _GEN_828; // @[FFT.scala 35:12]
  wire [31:0] _GEN_829; // @[FFT.scala 35:12]
  wire [31:0] _GEN_830; // @[FFT.scala 35:12]
  wire [31:0] _GEN_831; // @[FFT.scala 35:12]
  wire [31:0] _GEN_832; // @[FFT.scala 35:12]
  wire [31:0] _GEN_833; // @[FFT.scala 35:12]
  wire [31:0] _GEN_834; // @[FFT.scala 35:12]
  wire [31:0] _GEN_835; // @[FFT.scala 35:12]
  wire [31:0] _GEN_836; // @[FFT.scala 35:12]
  wire [31:0] _GEN_837; // @[FFT.scala 35:12]
  wire [31:0] _GEN_838; // @[FFT.scala 35:12]
  wire [31:0] _GEN_839; // @[FFT.scala 35:12]
  wire [31:0] _GEN_840; // @[FFT.scala 35:12]
  wire [31:0] _GEN_841; // @[FFT.scala 35:12]
  wire [31:0] _GEN_842; // @[FFT.scala 35:12]
  wire [31:0] _GEN_843; // @[FFT.scala 35:12]
  wire [31:0] _GEN_844; // @[FFT.scala 35:12]
  wire [31:0] _GEN_845; // @[FFT.scala 35:12]
  wire [31:0] _GEN_846; // @[FFT.scala 35:12]
  wire [31:0] _GEN_847; // @[FFT.scala 35:12]
  wire [31:0] _GEN_848; // @[FFT.scala 35:12]
  wire [31:0] _GEN_849; // @[FFT.scala 35:12]
  wire [31:0] _GEN_850; // @[FFT.scala 35:12]
  wire [31:0] _GEN_851; // @[FFT.scala 35:12]
  wire [31:0] _GEN_852; // @[FFT.scala 35:12]
  wire [31:0] _GEN_853; // @[FFT.scala 35:12]
  wire [31:0] _GEN_854; // @[FFT.scala 35:12]
  wire [31:0] _GEN_855; // @[FFT.scala 35:12]
  wire [31:0] _GEN_856; // @[FFT.scala 35:12]
  wire [31:0] _GEN_857; // @[FFT.scala 35:12]
  wire [31:0] _GEN_858; // @[FFT.scala 35:12]
  wire [31:0] _GEN_859; // @[FFT.scala 35:12]
  wire [31:0] _GEN_860; // @[FFT.scala 35:12]
  wire [31:0] _GEN_861; // @[FFT.scala 35:12]
  wire [31:0] _GEN_862; // @[FFT.scala 35:12]
  wire [31:0] _GEN_863; // @[FFT.scala 35:12]
  wire [31:0] _GEN_864; // @[FFT.scala 35:12]
  wire [31:0] _GEN_865; // @[FFT.scala 35:12]
  wire [31:0] _GEN_866; // @[FFT.scala 35:12]
  wire [31:0] _GEN_867; // @[FFT.scala 35:12]
  wire [31:0] _GEN_868; // @[FFT.scala 35:12]
  wire [31:0] _GEN_869; // @[FFT.scala 35:12]
  wire [31:0] _GEN_870; // @[FFT.scala 35:12]
  wire [31:0] _GEN_871; // @[FFT.scala 35:12]
  wire [31:0] _GEN_872; // @[FFT.scala 35:12]
  wire [31:0] _GEN_873; // @[FFT.scala 35:12]
  wire [31:0] _GEN_874; // @[FFT.scala 35:12]
  wire [31:0] _GEN_875; // @[FFT.scala 35:12]
  wire [31:0] _GEN_876; // @[FFT.scala 35:12]
  wire [31:0] _GEN_877; // @[FFT.scala 35:12]
  wire [31:0] _GEN_878; // @[FFT.scala 35:12]
  wire [31:0] _GEN_879; // @[FFT.scala 35:12]
  wire [31:0] _GEN_880; // @[FFT.scala 35:12]
  wire [31:0] _GEN_881; // @[FFT.scala 35:12]
  wire [31:0] _GEN_882; // @[FFT.scala 35:12]
  wire [31:0] _GEN_883; // @[FFT.scala 35:12]
  wire [31:0] _GEN_884; // @[FFT.scala 35:12]
  wire [31:0] _GEN_885; // @[FFT.scala 35:12]
  wire [31:0] _GEN_886; // @[FFT.scala 35:12]
  wire [31:0] _GEN_887; // @[FFT.scala 35:12]
  wire [31:0] _GEN_888; // @[FFT.scala 35:12]
  wire [31:0] _GEN_889; // @[FFT.scala 35:12]
  wire [31:0] _GEN_890; // @[FFT.scala 35:12]
  wire [31:0] _GEN_891; // @[FFT.scala 35:12]
  wire [31:0] _GEN_892; // @[FFT.scala 35:12]
  wire [31:0] _GEN_893; // @[FFT.scala 35:12]
  wire [31:0] _GEN_894; // @[FFT.scala 35:12]
  wire [31:0] _GEN_895; // @[FFT.scala 35:12]
  wire [31:0] _GEN_896; // @[FFT.scala 35:12]
  wire [31:0] _GEN_897; // @[FFT.scala 35:12]
  wire [31:0] _GEN_898; // @[FFT.scala 35:12]
  wire [31:0] _GEN_899; // @[FFT.scala 35:12]
  wire [31:0] _GEN_900; // @[FFT.scala 35:12]
  wire [31:0] _GEN_901; // @[FFT.scala 35:12]
  wire [31:0] _GEN_902; // @[FFT.scala 35:12]
  wire [31:0] _GEN_903; // @[FFT.scala 35:12]
  wire [31:0] _GEN_904; // @[FFT.scala 35:12]
  wire [31:0] _GEN_905; // @[FFT.scala 35:12]
  wire [31:0] _GEN_906; // @[FFT.scala 35:12]
  wire [31:0] _GEN_907; // @[FFT.scala 35:12]
  wire [31:0] _GEN_908; // @[FFT.scala 35:12]
  wire [31:0] _GEN_909; // @[FFT.scala 35:12]
  wire [31:0] _GEN_910; // @[FFT.scala 35:12]
  wire [31:0] _GEN_911; // @[FFT.scala 35:12]
  wire [31:0] _GEN_912; // @[FFT.scala 35:12]
  wire [31:0] _GEN_913; // @[FFT.scala 35:12]
  wire [31:0] _GEN_914; // @[FFT.scala 35:12]
  wire [31:0] _GEN_915; // @[FFT.scala 35:12]
  wire [31:0] _GEN_916; // @[FFT.scala 35:12]
  wire [31:0] _GEN_917; // @[FFT.scala 35:12]
  wire [31:0] _GEN_918; // @[FFT.scala 35:12]
  wire [31:0] _GEN_919; // @[FFT.scala 35:12]
  wire [31:0] _GEN_920; // @[FFT.scala 35:12]
  wire [31:0] _GEN_921; // @[FFT.scala 35:12]
  wire [31:0] _GEN_922; // @[FFT.scala 35:12]
  wire [31:0] _GEN_923; // @[FFT.scala 35:12]
  wire [31:0] _GEN_924; // @[FFT.scala 35:12]
  wire [31:0] _GEN_925; // @[FFT.scala 35:12]
  wire [31:0] _GEN_926; // @[FFT.scala 35:12]
  wire [31:0] _GEN_927; // @[FFT.scala 35:12]
  wire [31:0] _GEN_928; // @[FFT.scala 35:12]
  wire [31:0] _GEN_929; // @[FFT.scala 35:12]
  wire [31:0] _GEN_930; // @[FFT.scala 35:12]
  wire [31:0] _GEN_931; // @[FFT.scala 35:12]
  wire [31:0] _GEN_932; // @[FFT.scala 35:12]
  wire [31:0] _GEN_933; // @[FFT.scala 35:12]
  wire [31:0] _GEN_934; // @[FFT.scala 35:12]
  wire [31:0] _GEN_935; // @[FFT.scala 35:12]
  wire [31:0] _GEN_936; // @[FFT.scala 35:12]
  wire [31:0] _GEN_937; // @[FFT.scala 35:12]
  wire [31:0] _GEN_938; // @[FFT.scala 35:12]
  wire [31:0] _GEN_939; // @[FFT.scala 35:12]
  wire [31:0] _GEN_940; // @[FFT.scala 35:12]
  wire [31:0] _GEN_941; // @[FFT.scala 35:12]
  wire [31:0] _GEN_942; // @[FFT.scala 35:12]
  wire [31:0] _GEN_943; // @[FFT.scala 35:12]
  wire [31:0] _GEN_944; // @[FFT.scala 35:12]
  wire [31:0] _GEN_945; // @[FFT.scala 35:12]
  wire [31:0] _GEN_946; // @[FFT.scala 35:12]
  wire [31:0] _GEN_947; // @[FFT.scala 35:12]
  wire [31:0] _GEN_948; // @[FFT.scala 35:12]
  wire [31:0] _GEN_949; // @[FFT.scala 35:12]
  wire [31:0] _GEN_950; // @[FFT.scala 35:12]
  wire [31:0] _GEN_951; // @[FFT.scala 35:12]
  wire [31:0] _GEN_952; // @[FFT.scala 35:12]
  wire [31:0] _GEN_953; // @[FFT.scala 35:12]
  wire [31:0] _GEN_954; // @[FFT.scala 35:12]
  wire [31:0] _GEN_955; // @[FFT.scala 35:12]
  wire [31:0] _GEN_956; // @[FFT.scala 35:12]
  wire [31:0] _GEN_957; // @[FFT.scala 35:12]
  wire [31:0] _GEN_958; // @[FFT.scala 35:12]
  wire [31:0] _GEN_959; // @[FFT.scala 35:12]
  wire [31:0] _GEN_960; // @[FFT.scala 35:12]
  wire [31:0] _GEN_961; // @[FFT.scala 35:12]
  wire [31:0] _GEN_962; // @[FFT.scala 35:12]
  wire [31:0] _GEN_963; // @[FFT.scala 35:12]
  wire [31:0] _GEN_964; // @[FFT.scala 35:12]
  wire [31:0] _GEN_965; // @[FFT.scala 35:12]
  wire [31:0] _GEN_966; // @[FFT.scala 35:12]
  wire [31:0] _GEN_967; // @[FFT.scala 35:12]
  wire [31:0] _GEN_968; // @[FFT.scala 35:12]
  wire [31:0] _GEN_969; // @[FFT.scala 35:12]
  wire [31:0] _GEN_970; // @[FFT.scala 35:12]
  wire [31:0] _GEN_971; // @[FFT.scala 35:12]
  wire [31:0] _GEN_972; // @[FFT.scala 35:12]
  wire [31:0] _GEN_973; // @[FFT.scala 35:12]
  wire [31:0] _GEN_974; // @[FFT.scala 35:12]
  wire [31:0] _GEN_975; // @[FFT.scala 35:12]
  wire [31:0] _GEN_976; // @[FFT.scala 35:12]
  wire [31:0] _GEN_977; // @[FFT.scala 35:12]
  wire [31:0] _GEN_978; // @[FFT.scala 35:12]
  wire [31:0] _GEN_979; // @[FFT.scala 35:12]
  wire [31:0] _GEN_980; // @[FFT.scala 35:12]
  wire [31:0] _GEN_981; // @[FFT.scala 35:12]
  wire [31:0] _GEN_982; // @[FFT.scala 35:12]
  wire [31:0] _GEN_983; // @[FFT.scala 35:12]
  wire [31:0] _GEN_984; // @[FFT.scala 35:12]
  wire [31:0] _GEN_985; // @[FFT.scala 35:12]
  wire [31:0] _GEN_986; // @[FFT.scala 35:12]
  wire [31:0] _GEN_987; // @[FFT.scala 35:12]
  wire [31:0] _GEN_988; // @[FFT.scala 35:12]
  wire [31:0] _GEN_989; // @[FFT.scala 35:12]
  wire [31:0] _GEN_990; // @[FFT.scala 35:12]
  wire [31:0] _GEN_991; // @[FFT.scala 35:12]
  wire [31:0] _GEN_992; // @[FFT.scala 35:12]
  wire [31:0] _GEN_993; // @[FFT.scala 35:12]
  wire [31:0] _GEN_994; // @[FFT.scala 35:12]
  wire [31:0] _GEN_995; // @[FFT.scala 35:12]
  wire [31:0] _GEN_996; // @[FFT.scala 35:12]
  wire [31:0] _GEN_997; // @[FFT.scala 35:12]
  wire [31:0] _GEN_998; // @[FFT.scala 35:12]
  wire [31:0] _GEN_999; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1000; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1001; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1002; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1003; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1004; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1005; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1006; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1007; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1008; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1009; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1010; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1011; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1012; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1013; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1014; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1015; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1016; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1017; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1018; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1019; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1020; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1021; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1022; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1023; // @[FFT.scala 35:12]
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [31:0] _T_161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [31:0] _T_163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [31:0] _T_328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [31:0] _T_393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [31:0] _T_402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [31:0] _T_406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [31:0] _T_409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [31:0] _T_409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_521;
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_522;
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_523;
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_524;
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_525;
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_526;
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_527;
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_528;
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_529;
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_530;
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_531;
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_532;
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_533;
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_534;
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_535;
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_536;
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_537;
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_538;
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_539;
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_540;
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_541;
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_552;
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_553;
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_554;
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_557;
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_558;
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_559;
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_560;
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_561;
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_562;
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_563;
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_564;
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_565;
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_566;
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_567;
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_568;
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_569;
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_570;
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_571;
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_572;
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_573;
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_574;
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_575;
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_576;
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_577;
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_578;
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_579;
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_580;
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_581;
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_582;
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_583;
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_584;
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_585;
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_586;
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_587;
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_588;
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_589;
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_590;
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_591;
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_592;
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_593;
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_594;
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_595;
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_596;
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_597;
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_598;
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_599;
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_600;
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_601;
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_602;
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_603;
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_604;
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_605;
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_606;
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_607;
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_608;
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_609;
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_610;
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_611;
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_612;
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_613;
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_614;
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_615;
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_616;
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_617;
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_618;
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_619;
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_620;
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_621;
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_622;
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_623;
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_624;
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_625;
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_626;
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_627;
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_628;
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_629;
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_630;
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_631;
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_632;
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_633;
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_634;
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_635;
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_636;
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_637;
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_638;
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_639;
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_640;
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_641;
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_642;
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_643;
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_644;
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_645;
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_646;
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_647;
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_648;
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_649;
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_650;
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_651;
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_652;
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_653;
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_654;
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_655;
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_656;
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_657;
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_658;
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_659;
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_660;
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_661;
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_662;
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_663;
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_664;
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_665;
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_666;
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_667;
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_668;
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_669;
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_670;
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_671;
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_672;
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_673;
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_674;
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_675;
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_676;
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_677;
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_678;
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_679;
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_680;
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_681;
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_682;
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_683;
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_684;
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_685;
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_686;
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_687;
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_688;
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_689;
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_690;
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_691;
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_692;
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_693;
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_694;
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_695;
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_696;
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_697;
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_698;
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_699;
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_700;
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_701;
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_702;
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_703;
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_704;
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_705;
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_706;
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_707;
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_708;
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_709;
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_710;
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_711;
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_712;
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_713;
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_714;
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_715;
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_716;
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_717;
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_718;
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_719;
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_720;
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_721;
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_722;
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_723;
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_724;
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_725;
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_726;
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_727;
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_728;
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_729;
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_730;
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_731;
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_732;
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_733;
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_734;
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_735;
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_736;
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_737;
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_738;
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_739;
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_740;
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_741;
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_742;
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_743;
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_744;
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_745;
  reg [31:0] _T_533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_746;
  reg [31:0] _T_533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_747;
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_748;
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_749;
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_750;
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_751;
  reg [31:0] _T_536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_752;
  reg [31:0] _T_536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_753;
  reg [31:0] _T_537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_754;
  reg [31:0] _T_537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_755;
  reg [31:0] _T_538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_756;
  reg [31:0] _T_538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_757;
  reg [31:0] _T_539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_758;
  reg [31:0] _T_539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_759;
  reg [31:0] _T_540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_760;
  reg [31:0] _T_540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_761;
  reg [31:0] _T_541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_762;
  reg [31:0] _T_541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_763;
  reg [31:0] _T_542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_764;
  reg [31:0] _T_542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_765;
  reg [31:0] _T_543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_766;
  reg [31:0] _T_543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_767;
  reg [31:0] _T_544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_768;
  reg [31:0] _T_544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_769;
  reg [31:0] _T_545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  reg [31:0] _T_545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_771;
  reg [31:0] _T_546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_772;
  reg [31:0] _T_546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_773;
  reg [31:0] _T_547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  reg [31:0] _T_547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_781;
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_782;
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_783;
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_784;
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_785;
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_786;
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_787;
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_788;
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_789;
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_790;
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_791;
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_792;
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_793;
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_794;
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_795;
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_796;
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_797;
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_798;
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_799;
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_800;
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_801;
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_802;
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_803;
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_804;
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_805;
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_806;
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_807;
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_808;
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_809;
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_810;
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_811;
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_812;
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_813;
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_814;
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_815;
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_816;
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_817;
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_818;
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_819;
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_820;
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_821;
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_822;
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_823;
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_824;
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_825;
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_826;
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_827;
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_828;
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_829;
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_830;
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_831;
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_832;
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_833;
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_834;
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_835;
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_836;
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_837;
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_838;
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_839;
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_840;
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_841;
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_842;
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_843;
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_844;
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_845;
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_846;
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_847;
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_848;
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_849;
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_850;
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_851;
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_852;
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_853;
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_854;
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_855;
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_856;
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_857;
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_858;
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_859;
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_860;
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_861;
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_862;
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_863;
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_864;
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_865;
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_866;
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_867;
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_868;
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_869;
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_870;
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_871;
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_872;
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_873;
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_874;
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_875;
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_876;
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_877;
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_878;
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_879;
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_880;
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_881;
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_882;
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_883;
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_884;
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_885;
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_886;
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_887;
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_888;
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_889;
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_890;
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_891;
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_892;
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_893;
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_894;
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_895;
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_896;
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_897;
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_898;
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_899;
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_900;
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_901;
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_902;
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_903;
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_904;
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_905;
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_906;
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_907;
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_908;
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_909;
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_910;
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_911;
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_912;
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_913;
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_914;
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_915;
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_916;
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_917;
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_918;
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_919;
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_920;
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_921;
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_922;
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_923;
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_924;
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_925;
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_926;
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_927;
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_928;
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_929;
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_930;
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_931;
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_932;
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_933;
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_934;
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_935;
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_936;
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_937;
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_938;
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_939;
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_940;
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_941;
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_942;
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_943;
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_944;
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_945;
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_946;
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_947;
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_948;
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_949;
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_950;
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_951;
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_952;
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_953;
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_954;
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_955;
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_956;
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_957;
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_958;
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_959;
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_960;
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_961;
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_962;
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_963;
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_964;
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_965;
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_966;
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_967;
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_968;
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_969;
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_970;
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_971;
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_972;
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_973;
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_974;
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_975;
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_976;
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_977;
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_978;
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_979;
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_980;
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_981;
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_982;
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_983;
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_984;
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_985;
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_986;
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_987;
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_988;
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_989;
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_990;
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_991;
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_992;
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_993;
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_994;
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_995;
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_996;
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_997;
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_998;
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_999;
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1000;
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1001;
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1002;
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1003;
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1004;
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1005;
  reg [31:0] _T_663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1006;
  reg [31:0] _T_663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1007;
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1008;
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1009;
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1010;
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1011;
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1012;
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1013;
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1014;
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1015;
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1016;
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1017;
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1018;
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1019;
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1020;
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1021;
  reg [31:0] _T_671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1022;
  reg [31:0] _T_671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1023;
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1024;
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1025;
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1026;
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1027;
  reg [31:0] _T_676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1028;
  reg [31:0] _T_676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1029;
  reg [31:0] _T_677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1030;
  reg [31:0] _T_677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1031;
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1032;
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1033;
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1034;
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1035;
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1036;
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1037;
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1038;
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1039;
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1040;
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1041;
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1042;
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1043;
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1044;
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1045;
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1046;
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1047;
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1048;
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1049;
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1050;
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1051;
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1052;
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1053;
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1054;
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1055;
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1056;
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1057;
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1058;
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1059;
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1060;
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1061;
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1062;
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1063;
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1064;
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1065;
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1066;
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1067;
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1068;
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1069;
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1070;
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1071;
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1072;
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1073;
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1074;
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1075;
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1076;
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1077;
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1078;
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1079;
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1080;
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1081;
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1082;
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1083;
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1084;
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1085;
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1086;
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1087;
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1088;
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1089;
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1090;
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1091;
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1092;
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1093;
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1094;
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1095;
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1096;
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1097;
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1098;
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1099;
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1100;
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1101;
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1102;
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1103;
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1104;
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1105;
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1106;
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1107;
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1108;
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1109;
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1110;
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1111;
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1112;
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1113;
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1114;
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1115;
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1116;
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1117;
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1118;
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1119;
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1120;
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1121;
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1122;
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1123;
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1124;
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1125;
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1126;
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1127;
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1128;
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1129;
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1130;
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1131;
  reg [31:0] _T_728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1132;
  reg [31:0] _T_728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1133;
  reg [31:0] _T_729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1134;
  reg [31:0] _T_729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1135;
  reg [31:0] _T_730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1136;
  reg [31:0] _T_730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1137;
  reg [31:0] _T_731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1138;
  reg [31:0] _T_731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1139;
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1140;
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1141;
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1142;
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1143;
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1144;
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1145;
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1146;
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1147;
  reg [31:0] _T_736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1148;
  reg [31:0] _T_736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1149;
  reg [31:0] _T_737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1150;
  reg [31:0] _T_737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1151;
  reg [31:0] _T_738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1152;
  reg [31:0] _T_738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1153;
  reg [31:0] _T_739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1154;
  reg [31:0] _T_739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1155;
  reg [31:0] _T_740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1156;
  reg [31:0] _T_740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1157;
  reg [31:0] _T_741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1158;
  reg [31:0] _T_741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1159;
  reg [31:0] _T_742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1160;
  reg [31:0] _T_742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1161;
  reg [31:0] _T_743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1162;
  reg [31:0] _T_743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1163;
  reg [31:0] _T_744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1164;
  reg [31:0] _T_744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1165;
  reg [31:0] _T_745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1166;
  reg [31:0] _T_745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1167;
  reg [31:0] _T_746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1168;
  reg [31:0] _T_746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1169;
  reg [31:0] _T_747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1170;
  reg [31:0] _T_747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1171;
  reg [31:0] _T_748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1172;
  reg [31:0] _T_748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1173;
  reg [31:0] _T_749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1174;
  reg [31:0] _T_749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1175;
  reg [31:0] _T_750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1176;
  reg [31:0] _T_750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1177;
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1178;
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1179;
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1180;
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1181;
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1182;
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1183;
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1184;
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1185;
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1186;
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1187;
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1188;
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1189;
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1190;
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1191;
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1192;
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1193;
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1194;
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1195;
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1196;
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1197;
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1198;
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1199;
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1200;
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1201;
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1202;
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1203;
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1204;
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1205;
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1206;
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1207;
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1208;
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1209;
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1210;
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1211;
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1212;
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1213;
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1214;
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1215;
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1216;
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1217;
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1218;
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1219;
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1220;
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1221;
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1222;
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1223;
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1224;
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1225;
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1226;
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1227;
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1228;
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1229;
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1230;
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1231;
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1232;
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1233;
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1234;
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1235;
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1236;
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1237;
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1238;
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1239;
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1240;
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1241;
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1242;
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1243;
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1244;
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1245;
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1246;
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1247;
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1248;
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1249;
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1250;
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1251;
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1252;
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1253;
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1254;
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1255;
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1256;
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1257;
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1258;
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1259;
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1260;
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1261;
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1262;
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1263;
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1264;
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1265;
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1266;
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1267;
  reg [31:0] _T_796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1268;
  reg [31:0] _T_796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1269;
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1270;
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1271;
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1272;
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1273;
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1274;
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1275;
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1276;
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1277;
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1278;
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1279;
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1280;
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1281;
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1282;
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1283;
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1284;
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1285;
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1286;
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1287;
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1288;
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1289;
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1290;
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1291;
  reg [31:0] _T_808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1292;
  reg [31:0] _T_808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1293;
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1294;
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1295;
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1296;
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1297;
  reg [31:0] _T_811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1298;
  reg [31:0] _T_811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1299;
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1300;
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1301;
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1302;
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1303;
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1304;
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1305;
  reg [31:0] _T_815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1306;
  reg [31:0] _T_815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1307;
  reg [31:0] _T_816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1308;
  reg [31:0] _T_816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1309;
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1310;
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1311;
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1312;
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1313;
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1314;
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1315;
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1316;
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1317;
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1318;
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1319;
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1320;
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1321;
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1322;
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1323;
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1324;
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1325;
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1326;
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1327;
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1328;
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1329;
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1330;
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1331;
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1332;
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1333;
  reg [31:0] _T_829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1334;
  reg [31:0] _T_829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1335;
  reg [31:0] _T_830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1336;
  reg [31:0] _T_830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1337;
  reg [31:0] _T_831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1338;
  reg [31:0] _T_831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1339;
  reg [31:0] _T_832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1340;
  reg [31:0] _T_832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1341;
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1342;
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1343;
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1344;
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1345;
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1346;
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1347;
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1348;
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1349;
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1350;
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1351;
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1352;
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1353;
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1354;
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1355;
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1356;
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1357;
  reg [31:0] _T_841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1358;
  reg [31:0] _T_841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1359;
  reg [31:0] _T_842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1360;
  reg [31:0] _T_842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1361;
  reg [31:0] _T_843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1362;
  reg [31:0] _T_843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1363;
  reg [31:0] _T_844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1364;
  reg [31:0] _T_844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1365;
  reg [31:0] _T_845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1366;
  reg [31:0] _T_845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1367;
  reg [31:0] _T_846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1368;
  reg [31:0] _T_846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1369;
  reg [31:0] _T_847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1370;
  reg [31:0] _T_847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1371;
  reg [31:0] _T_848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1372;
  reg [31:0] _T_848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1373;
  reg [31:0] _T_849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1374;
  reg [31:0] _T_849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1375;
  reg [31:0] _T_850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1376;
  reg [31:0] _T_850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1377;
  reg [31:0] _T_851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1378;
  reg [31:0] _T_851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1379;
  reg [31:0] _T_852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1380;
  reg [31:0] _T_852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1381;
  reg [31:0] _T_853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1382;
  reg [31:0] _T_853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1383;
  reg [31:0] _T_854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1384;
  reg [31:0] _T_854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1385;
  reg [31:0] _T_855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1386;
  reg [31:0] _T_855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1387;
  reg [31:0] _T_856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1388;
  reg [31:0] _T_856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1389;
  reg [31:0] _T_857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1390;
  reg [31:0] _T_857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1391;
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1392;
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1393;
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1394;
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1395;
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1396;
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1397;
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1398;
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1399;
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1400;
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1401;
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1402;
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1403;
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1404;
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1405;
  reg [31:0] _T_865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1406;
  reg [31:0] _T_865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1407;
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1408;
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1409;
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1410;
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1411;
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1412;
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1413;
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1414;
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1415;
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1416;
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1417;
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1418;
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1419;
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1420;
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1421;
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1422;
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1423;
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1424;
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1425;
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1426;
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1427;
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1428;
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1429;
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1430;
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1431;
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1432;
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1433;
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1434;
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1435;
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1436;
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1437;
  reg [31:0] _T_881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1438;
  reg [31:0] _T_881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1439;
  reg [31:0] _T_882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1440;
  reg [31:0] _T_882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1441;
  reg [31:0] _T_883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1442;
  reg [31:0] _T_883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1443;
  reg [31:0] _T_884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1444;
  reg [31:0] _T_884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1445;
  reg [31:0] _T_885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1446;
  reg [31:0] _T_885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1447;
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1448;
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1449;
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1450;
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1451;
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1452;
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1453;
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1454;
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1455;
  reg [31:0] _T_890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1456;
  reg [31:0] _T_890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1457;
  reg [31:0] _T_891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1458;
  reg [31:0] _T_891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1459;
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1460;
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1461;
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1462;
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1463;
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1464;
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1465;
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1466;
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1467;
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1468;
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1469;
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1470;
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1471;
  reg [31:0] _T_898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1472;
  reg [31:0] _T_898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1473;
  reg [31:0] _T_899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1474;
  reg [31:0] _T_899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1475;
  reg [31:0] _T_900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1476;
  reg [31:0] _T_900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1477;
  reg [31:0] _T_901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1478;
  reg [31:0] _T_901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1479;
  reg [31:0] _T_902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1480;
  reg [31:0] _T_902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1481;
  reg [31:0] _T_903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1482;
  reg [31:0] _T_903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1483;
  reg [31:0] _T_904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1484;
  reg [31:0] _T_904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1485;
  reg [31:0] _T_905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1486;
  reg [31:0] _T_905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1487;
  reg [31:0] _T_906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1488;
  reg [31:0] _T_906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1489;
  reg [31:0] _T_907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1490;
  reg [31:0] _T_907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1491;
  reg [31:0] _T_908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1492;
  reg [31:0] _T_908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1493;
  reg [31:0] _T_909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1494;
  reg [31:0] _T_909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1495;
  reg [31:0] _T_910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1496;
  reg [31:0] _T_910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1497;
  reg [31:0] _T_911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1498;
  reg [31:0] _T_911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1499;
  reg [31:0] _T_912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1500;
  reg [31:0] _T_912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1501;
  reg [31:0] _T_913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1502;
  reg [31:0] _T_913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1503;
  reg [31:0] _T_914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1504;
  reg [31:0] _T_914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1505;
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1506;
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1507;
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1508;
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1509;
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1510;
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1511;
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1512;
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1513;
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1514;
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1515;
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1516;
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1517;
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1518;
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1519;
  reg [31:0] _T_922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1520;
  reg [31:0] _T_922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1521;
  reg [31:0] _T_923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1522;
  reg [31:0] _T_923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1523;
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1524;
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1525;
  reg [31:0] _T_925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1526;
  reg [31:0] _T_925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1527;
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1528;
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1529;
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1530;
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1531;
  reg [31:0] _T_928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1532;
  reg [31:0] _T_928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1533;
  reg [31:0] _T_929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1534;
  reg [31:0] _T_929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1535;
  reg [31:0] _T_930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1536;
  reg [31:0] _T_930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1537;
  wire [31:0] _GEN_2562; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2563; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2564; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2565; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2566; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2567; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2568; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2569; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2570; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2571; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2572; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2573; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2574; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2575; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2576; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2577; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2578; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2579; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2580; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2581; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2582; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2583; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2584; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2585; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2586; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2587; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2588; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2589; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2590; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2591; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2592; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2593; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2594; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2595; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2596; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2597; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2598; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2599; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2600; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2601; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2602; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2603; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2604; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2605; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2606; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2607; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2608; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2609; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2610; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2611; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2612; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2613; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2614; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2615; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2616; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2617; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2618; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2619; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2620; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2621; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2622; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2623; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2624; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2625; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2626; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2627; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2628; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2629; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2630; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2631; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2632; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2633; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2634; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2635; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2636; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2637; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2638; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2639; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2640; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2641; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2642; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2643; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2644; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2645; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2646; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2647; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2648; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2649; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2650; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2651; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2652; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2653; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2654; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2655; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2656; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2657; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2658; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2659; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2660; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2661; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2662; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2663; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2664; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2665; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2666; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2667; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2668; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2669; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2670; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2671; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2672; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2673; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2674; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2675; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2676; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2677; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2678; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2679; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2680; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2681; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2682; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2683; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2684; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2685; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2686; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2687; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2688; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2689; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2690; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2691; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2692; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2693; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2694; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2695; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2696; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2697; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2698; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2699; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2700; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2701; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2702; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2703; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2704; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2705; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2706; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2707; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2708; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2709; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2710; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2711; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2712; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2713; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2714; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2715; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2716; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2717; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2718; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2719; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2720; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2721; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2722; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2723; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2724; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2725; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2726; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2727; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2728; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2729; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2730; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2731; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2732; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2733; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2734; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2735; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2736; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2737; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2738; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2739; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2740; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2741; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2742; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2743; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2744; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2745; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2746; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2747; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2748; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2749; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2750; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2751; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2752; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2753; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2754; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2755; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2756; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2757; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2758; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2759; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2760; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2761; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2762; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2763; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2764; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2765; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2766; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2767; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2768; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2769; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2770; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2771; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2772; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2773; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2774; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2775; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2776; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2777; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2778; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2779; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2780; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2781; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2782; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2783; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2784; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2785; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2786; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2787; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2788; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2789; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2790; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2791; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2792; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2793; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2794; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2795; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2796; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2797; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2798; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2799; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2800; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2801; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2802; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2803; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2804; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2805; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2806; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2807; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2808; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2809; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2810; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2811; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2812; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2813; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2814; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2815; // @[FFT.scala 34:12]
  wire [31:0] _GEN_2818; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2819; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2820; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2821; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2822; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2823; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2824; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2825; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2826; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2827; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2828; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2829; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2830; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2831; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2832; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2833; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2834; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2835; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2836; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2837; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2838; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2839; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2840; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2841; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2842; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2843; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2844; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2845; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2846; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2847; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2848; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2849; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2850; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2851; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2852; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2853; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2854; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2855; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2856; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2857; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2858; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2859; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2860; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2861; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2862; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2863; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2864; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2865; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2866; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2867; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2868; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2869; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2870; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2871; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2872; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2873; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2874; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2875; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2876; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2877; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2878; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2879; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2880; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2881; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2882; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2883; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2884; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2885; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2886; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2887; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2888; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2889; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2890; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2891; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2892; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2893; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2894; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2895; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2896; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2897; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2898; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2899; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2900; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2901; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2902; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2903; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2904; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2905; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2906; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2907; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2908; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2909; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2910; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2911; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2912; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2913; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2914; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2915; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2916; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2917; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2918; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2919; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2920; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2921; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2922; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2923; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2924; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2925; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2926; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2927; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2928; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2929; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2930; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2931; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2932; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2933; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2934; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2935; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2936; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2937; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2938; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2939; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2940; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2941; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2942; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2943; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2944; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2945; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2946; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2947; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2948; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2949; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2950; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2951; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2952; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2953; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2954; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2955; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2956; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2957; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2958; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2959; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2960; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2961; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2962; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2963; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2964; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2965; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2966; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2967; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2968; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2969; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2970; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2971; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2972; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2973; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2974; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2975; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2976; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2977; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2978; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2979; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2980; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2981; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2982; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2983; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2984; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2985; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2986; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2987; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2988; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2989; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2990; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2991; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2992; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2993; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2994; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2995; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2996; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2997; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2998; // @[FFT.scala 35:12]
  wire [31:0] _GEN_2999; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3000; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3001; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3002; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3003; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3004; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3005; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3006; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3007; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3008; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3009; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3010; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3011; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3012; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3013; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3014; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3015; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3016; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3017; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3018; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3019; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3020; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3021; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3022; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3023; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3024; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3025; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3026; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3027; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3028; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3029; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3030; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3031; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3032; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3033; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3034; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3035; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3036; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3037; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3038; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3039; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3040; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3041; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3042; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3043; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3044; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3045; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3046; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3047; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3048; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3049; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3050; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3051; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3052; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3053; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3054; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3055; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3056; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3057; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3058; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3059; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3060; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3061; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3062; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3063; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3064; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3065; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3066; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3067; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3068; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3069; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3070; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3071; // @[FFT.scala 35:12]
  reg [31:0] _T_936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1538;
  reg [31:0] _T_936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1539;
  reg [31:0] _T_937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1540;
  reg [31:0] _T_937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1541;
  reg [31:0] _T_938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1542;
  reg [31:0] _T_938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1543;
  reg [31:0] _T_939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1544;
  reg [31:0] _T_939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1545;
  reg [31:0] _T_940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1546;
  reg [31:0] _T_940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1547;
  reg [31:0] _T_941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1548;
  reg [31:0] _T_941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1549;
  reg [31:0] _T_942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1550;
  reg [31:0] _T_942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1551;
  reg [31:0] _T_943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1552;
  reg [31:0] _T_943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1553;
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1554;
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1555;
  reg [31:0] _T_945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1556;
  reg [31:0] _T_945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1557;
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1558;
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1559;
  reg [31:0] _T_947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1560;
  reg [31:0] _T_947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1561;
  reg [31:0] _T_948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1562;
  reg [31:0] _T_948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1563;
  reg [31:0] _T_949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1564;
  reg [31:0] _T_949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1565;
  reg [31:0] _T_950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1566;
  reg [31:0] _T_950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1567;
  reg [31:0] _T_951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1568;
  reg [31:0] _T_951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1569;
  reg [31:0] _T_952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1570;
  reg [31:0] _T_952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1571;
  reg [31:0] _T_953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1572;
  reg [31:0] _T_953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1573;
  reg [31:0] _T_954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1574;
  reg [31:0] _T_954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1575;
  reg [31:0] _T_955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1576;
  reg [31:0] _T_955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1577;
  reg [31:0] _T_956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1578;
  reg [31:0] _T_956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1579;
  reg [31:0] _T_957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1580;
  reg [31:0] _T_957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1581;
  reg [31:0] _T_958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1582;
  reg [31:0] _T_958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1583;
  reg [31:0] _T_959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1584;
  reg [31:0] _T_959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1585;
  reg [31:0] _T_960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1586;
  reg [31:0] _T_960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1587;
  reg [31:0] _T_961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1588;
  reg [31:0] _T_961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1589;
  reg [31:0] _T_962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1590;
  reg [31:0] _T_962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1591;
  reg [31:0] _T_963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1592;
  reg [31:0] _T_963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1593;
  reg [31:0] _T_964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1594;
  reg [31:0] _T_964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1595;
  reg [31:0] _T_965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1596;
  reg [31:0] _T_965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1597;
  reg [31:0] _T_966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1598;
  reg [31:0] _T_966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1599;
  reg [31:0] _T_967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1600;
  reg [31:0] _T_967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1601;
  reg [31:0] _T_968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1602;
  reg [31:0] _T_968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1603;
  reg [31:0] _T_969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1604;
  reg [31:0] _T_969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1605;
  reg [31:0] _T_970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1606;
  reg [31:0] _T_970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1607;
  reg [31:0] _T_971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1608;
  reg [31:0] _T_971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1609;
  reg [31:0] _T_972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1610;
  reg [31:0] _T_972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1611;
  reg [31:0] _T_973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1612;
  reg [31:0] _T_973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1613;
  reg [31:0] _T_974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1614;
  reg [31:0] _T_974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1615;
  reg [31:0] _T_975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1616;
  reg [31:0] _T_975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1617;
  reg [31:0] _T_976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1618;
  reg [31:0] _T_976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1619;
  reg [31:0] _T_977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1620;
  reg [31:0] _T_977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1621;
  reg [31:0] _T_978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1622;
  reg [31:0] _T_978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1623;
  reg [31:0] _T_979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1624;
  reg [31:0] _T_979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1625;
  reg [31:0] _T_980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1626;
  reg [31:0] _T_980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1627;
  reg [31:0] _T_981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1628;
  reg [31:0] _T_981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1629;
  reg [31:0] _T_982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1630;
  reg [31:0] _T_982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1631;
  reg [31:0] _T_983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1632;
  reg [31:0] _T_983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1633;
  reg [31:0] _T_984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1634;
  reg [31:0] _T_984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1635;
  reg [31:0] _T_985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1636;
  reg [31:0] _T_985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1637;
  reg [31:0] _T_986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1638;
  reg [31:0] _T_986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1639;
  reg [31:0] _T_987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1640;
  reg [31:0] _T_987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1641;
  reg [31:0] _T_988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1642;
  reg [31:0] _T_988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1643;
  reg [31:0] _T_989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1644;
  reg [31:0] _T_989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1645;
  reg [31:0] _T_990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1646;
  reg [31:0] _T_990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1647;
  reg [31:0] _T_991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1648;
  reg [31:0] _T_991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1649;
  reg [31:0] _T_992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1650;
  reg [31:0] _T_992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1651;
  reg [31:0] _T_993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1652;
  reg [31:0] _T_993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1653;
  reg [31:0] _T_994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1654;
  reg [31:0] _T_994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1655;
  reg [31:0] _T_995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1656;
  reg [31:0] _T_995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1657;
  reg [31:0] _T_996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1658;
  reg [31:0] _T_996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1659;
  reg [31:0] _T_997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1660;
  reg [31:0] _T_997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1661;
  reg [31:0] _T_998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1662;
  reg [31:0] _T_998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1663;
  reg [31:0] _T_999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1664;
  reg [31:0] _T_999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1665;
  reg [31:0] _T_1000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1666;
  reg [31:0] _T_1000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1667;
  reg [31:0] _T_1001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1668;
  reg [31:0] _T_1001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1669;
  reg [31:0] _T_1002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1670;
  reg [31:0] _T_1002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1671;
  reg [31:0] _T_1003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1672;
  reg [31:0] _T_1003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1673;
  reg [31:0] _T_1004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1674;
  reg [31:0] _T_1004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1675;
  reg [31:0] _T_1005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1676;
  reg [31:0] _T_1005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1677;
  reg [31:0] _T_1006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1678;
  reg [31:0] _T_1006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1679;
  reg [31:0] _T_1007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1680;
  reg [31:0] _T_1007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1681;
  reg [31:0] _T_1008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1682;
  reg [31:0] _T_1008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1683;
  reg [31:0] _T_1009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1684;
  reg [31:0] _T_1009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1685;
  reg [31:0] _T_1010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1686;
  reg [31:0] _T_1010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1687;
  reg [31:0] _T_1011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1688;
  reg [31:0] _T_1011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1689;
  reg [31:0] _T_1012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1690;
  reg [31:0] _T_1012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1691;
  reg [31:0] _T_1013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1692;
  reg [31:0] _T_1013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1693;
  reg [31:0] _T_1014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1694;
  reg [31:0] _T_1014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1695;
  reg [31:0] _T_1015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1696;
  reg [31:0] _T_1015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1697;
  reg [31:0] _T_1016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1698;
  reg [31:0] _T_1016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1699;
  reg [31:0] _T_1017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1700;
  reg [31:0] _T_1017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1701;
  reg [31:0] _T_1018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1702;
  reg [31:0] _T_1018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1703;
  reg [31:0] _T_1019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1704;
  reg [31:0] _T_1019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1705;
  reg [31:0] _T_1020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1706;
  reg [31:0] _T_1020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1707;
  reg [31:0] _T_1021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1708;
  reg [31:0] _T_1021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1709;
  reg [31:0] _T_1022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1710;
  reg [31:0] _T_1022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1711;
  reg [31:0] _T_1023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1712;
  reg [31:0] _T_1023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1713;
  reg [31:0] _T_1024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1714;
  reg [31:0] _T_1024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1715;
  reg [31:0] _T_1025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1716;
  reg [31:0] _T_1025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1717;
  reg [31:0] _T_1026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1718;
  reg [31:0] _T_1026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1719;
  reg [31:0] _T_1027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1720;
  reg [31:0] _T_1027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1721;
  reg [31:0] _T_1028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1722;
  reg [31:0] _T_1028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1723;
  reg [31:0] _T_1029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1724;
  reg [31:0] _T_1029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1725;
  reg [31:0] _T_1030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1726;
  reg [31:0] _T_1030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1727;
  reg [31:0] _T_1031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1728;
  reg [31:0] _T_1031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1729;
  reg [31:0] _T_1032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1730;
  reg [31:0] _T_1032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1731;
  reg [31:0] _T_1033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1732;
  reg [31:0] _T_1033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1733;
  reg [31:0] _T_1034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1734;
  reg [31:0] _T_1034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1735;
  reg [31:0] _T_1035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1736;
  reg [31:0] _T_1035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1737;
  reg [31:0] _T_1036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1738;
  reg [31:0] _T_1036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1739;
  reg [31:0] _T_1037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1740;
  reg [31:0] _T_1037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1741;
  reg [31:0] _T_1038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1742;
  reg [31:0] _T_1038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1743;
  reg [31:0] _T_1039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1744;
  reg [31:0] _T_1039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1745;
  reg [31:0] _T_1040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1746;
  reg [31:0] _T_1040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1747;
  reg [31:0] _T_1041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1748;
  reg [31:0] _T_1041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1749;
  reg [31:0] _T_1042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1750;
  reg [31:0] _T_1042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1751;
  reg [31:0] _T_1043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1752;
  reg [31:0] _T_1043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1753;
  reg [31:0] _T_1044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1754;
  reg [31:0] _T_1044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1755;
  reg [31:0] _T_1045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1756;
  reg [31:0] _T_1045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1757;
  reg [31:0] _T_1046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1758;
  reg [31:0] _T_1046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1759;
  reg [31:0] _T_1047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1760;
  reg [31:0] _T_1047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1761;
  reg [31:0] _T_1048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1762;
  reg [31:0] _T_1048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1763;
  reg [31:0] _T_1049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1764;
  reg [31:0] _T_1049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1765;
  reg [31:0] _T_1050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1766;
  reg [31:0] _T_1050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1767;
  reg [31:0] _T_1051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1768;
  reg [31:0] _T_1051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1769;
  reg [31:0] _T_1052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1770;
  reg [31:0] _T_1052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1771;
  reg [31:0] _T_1053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1772;
  reg [31:0] _T_1053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1773;
  reg [31:0] _T_1054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1774;
  reg [31:0] _T_1054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1775;
  reg [31:0] _T_1055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1776;
  reg [31:0] _T_1055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1777;
  reg [31:0] _T_1056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1778;
  reg [31:0] _T_1056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1779;
  reg [31:0] _T_1057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1780;
  reg [31:0] _T_1057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1781;
  reg [31:0] _T_1058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1782;
  reg [31:0] _T_1058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1783;
  reg [31:0] _T_1059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1784;
  reg [31:0] _T_1059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1785;
  reg [31:0] _T_1060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1786;
  reg [31:0] _T_1060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1787;
  reg [31:0] _T_1061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1788;
  reg [31:0] _T_1061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1789;
  reg [31:0] _T_1062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1790;
  reg [31:0] _T_1062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1791;
  reg [31:0] _T_1063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1792;
  reg [31:0] _T_1063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1793;
  reg [31:0] _T_1064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1794;
  reg [31:0] _T_1064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1795;
  reg [31:0] _T_1065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1796;
  reg [31:0] _T_1065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1797;
  reg [31:0] _T_1066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1798;
  reg [31:0] _T_1066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1799;
  reg [31:0] _T_1067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1800;
  reg [31:0] _T_1067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1801;
  reg [31:0] _T_1068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1802;
  reg [31:0] _T_1068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1803;
  reg [31:0] _T_1069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1804;
  reg [31:0] _T_1069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1805;
  reg [31:0] _T_1070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1806;
  reg [31:0] _T_1070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1807;
  reg [31:0] _T_1071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1808;
  reg [31:0] _T_1071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1809;
  reg [31:0] _T_1072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1810;
  reg [31:0] _T_1072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1811;
  reg [31:0] _T_1073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1812;
  reg [31:0] _T_1073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1813;
  reg [31:0] _T_1074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1814;
  reg [31:0] _T_1074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1815;
  reg [31:0] _T_1075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1816;
  reg [31:0] _T_1075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1817;
  reg [31:0] _T_1076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1818;
  reg [31:0] _T_1076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1819;
  reg [31:0] _T_1077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1820;
  reg [31:0] _T_1077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1821;
  reg [31:0] _T_1078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1822;
  reg [31:0] _T_1078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1823;
  reg [31:0] _T_1079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1824;
  reg [31:0] _T_1079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1825;
  reg [31:0] _T_1080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1826;
  reg [31:0] _T_1080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1827;
  reg [31:0] _T_1081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1828;
  reg [31:0] _T_1081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1829;
  reg [31:0] _T_1082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1830;
  reg [31:0] _T_1082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1831;
  reg [31:0] _T_1083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1832;
  reg [31:0] _T_1083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1833;
  reg [31:0] _T_1084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1834;
  reg [31:0] _T_1084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1835;
  reg [31:0] _T_1085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1836;
  reg [31:0] _T_1085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1837;
  reg [31:0] _T_1086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1838;
  reg [31:0] _T_1086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1839;
  reg [31:0] _T_1087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1840;
  reg [31:0] _T_1087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1841;
  reg [31:0] _T_1088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1842;
  reg [31:0] _T_1088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1843;
  reg [31:0] _T_1089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1844;
  reg [31:0] _T_1089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1845;
  reg [31:0] _T_1090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1846;
  reg [31:0] _T_1090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1847;
  reg [31:0] _T_1091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1848;
  reg [31:0] _T_1091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1849;
  reg [31:0] _T_1092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1850;
  reg [31:0] _T_1092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1851;
  reg [31:0] _T_1093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1852;
  reg [31:0] _T_1093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1853;
  reg [31:0] _T_1094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1854;
  reg [31:0] _T_1094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1855;
  reg [31:0] _T_1095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1856;
  reg [31:0] _T_1095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1857;
  reg [31:0] _T_1096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1858;
  reg [31:0] _T_1096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1859;
  reg [31:0] _T_1097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1860;
  reg [31:0] _T_1097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1861;
  reg [31:0] _T_1098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1862;
  reg [31:0] _T_1098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1863;
  reg [31:0] _T_1099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1864;
  reg [31:0] _T_1099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1865;
  reg [31:0] _T_1100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1866;
  reg [31:0] _T_1100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1867;
  reg [31:0] _T_1101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1868;
  reg [31:0] _T_1101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1869;
  reg [31:0] _T_1102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1870;
  reg [31:0] _T_1102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1871;
  reg [31:0] _T_1103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1872;
  reg [31:0] _T_1103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1873;
  reg [31:0] _T_1104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1874;
  reg [31:0] _T_1104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1875;
  reg [31:0] _T_1105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1876;
  reg [31:0] _T_1105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1877;
  reg [31:0] _T_1106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1878;
  reg [31:0] _T_1106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1879;
  reg [31:0] _T_1107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1880;
  reg [31:0] _T_1107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1881;
  reg [31:0] _T_1108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1882;
  reg [31:0] _T_1108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1883;
  reg [31:0] _T_1109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1884;
  reg [31:0] _T_1109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1885;
  reg [31:0] _T_1110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1886;
  reg [31:0] _T_1110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1887;
  reg [31:0] _T_1111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1888;
  reg [31:0] _T_1111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1889;
  reg [31:0] _T_1112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1890;
  reg [31:0] _T_1112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1891;
  reg [31:0] _T_1113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1892;
  reg [31:0] _T_1113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1893;
  reg [31:0] _T_1114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1894;
  reg [31:0] _T_1114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1895;
  reg [31:0] _T_1115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1896;
  reg [31:0] _T_1115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1897;
  reg [31:0] _T_1116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1898;
  reg [31:0] _T_1116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1899;
  reg [31:0] _T_1117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1900;
  reg [31:0] _T_1117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1901;
  reg [31:0] _T_1118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1902;
  reg [31:0] _T_1118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1903;
  reg [31:0] _T_1119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1904;
  reg [31:0] _T_1119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1905;
  reg [31:0] _T_1120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1906;
  reg [31:0] _T_1120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1907;
  reg [31:0] _T_1121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1908;
  reg [31:0] _T_1121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1909;
  reg [31:0] _T_1122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1910;
  reg [31:0] _T_1122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1911;
  reg [31:0] _T_1123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1912;
  reg [31:0] _T_1123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1913;
  reg [31:0] _T_1124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1914;
  reg [31:0] _T_1124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1915;
  reg [31:0] _T_1125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1916;
  reg [31:0] _T_1125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1917;
  reg [31:0] _T_1126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1918;
  reg [31:0] _T_1126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1919;
  reg [31:0] _T_1127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1920;
  reg [31:0] _T_1127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1921;
  reg [31:0] _T_1128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1922;
  reg [31:0] _T_1128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1923;
  reg [31:0] _T_1129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1924;
  reg [31:0] _T_1129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1925;
  reg [31:0] _T_1130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1926;
  reg [31:0] _T_1130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1927;
  reg [31:0] _T_1131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1928;
  reg [31:0] _T_1131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1929;
  reg [31:0] _T_1132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1930;
  reg [31:0] _T_1132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1931;
  reg [31:0] _T_1133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1932;
  reg [31:0] _T_1133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1933;
  reg [31:0] _T_1134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1934;
  reg [31:0] _T_1134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1935;
  reg [31:0] _T_1135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1936;
  reg [31:0] _T_1135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1937;
  reg [31:0] _T_1136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1938;
  reg [31:0] _T_1136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1939;
  reg [31:0] _T_1137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1940;
  reg [31:0] _T_1137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1941;
  reg [31:0] _T_1138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1942;
  reg [31:0] _T_1138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1943;
  reg [31:0] _T_1139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1944;
  reg [31:0] _T_1139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1945;
  reg [31:0] _T_1140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1946;
  reg [31:0] _T_1140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1947;
  reg [31:0] _T_1141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1948;
  reg [31:0] _T_1141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1949;
  reg [31:0] _T_1142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1950;
  reg [31:0] _T_1142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1951;
  reg [31:0] _T_1143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1952;
  reg [31:0] _T_1143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1953;
  reg [31:0] _T_1144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1954;
  reg [31:0] _T_1144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1955;
  reg [31:0] _T_1145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1956;
  reg [31:0] _T_1145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1957;
  reg [31:0] _T_1146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1958;
  reg [31:0] _T_1146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1959;
  reg [31:0] _T_1147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1960;
  reg [31:0] _T_1147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1961;
  reg [31:0] _T_1148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1962;
  reg [31:0] _T_1148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1963;
  reg [31:0] _T_1149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1964;
  reg [31:0] _T_1149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1965;
  reg [31:0] _T_1150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1966;
  reg [31:0] _T_1150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1967;
  reg [31:0] _T_1151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1968;
  reg [31:0] _T_1151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1969;
  reg [31:0] _T_1152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1970;
  reg [31:0] _T_1152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1971;
  reg [31:0] _T_1153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1972;
  reg [31:0] _T_1153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1973;
  reg [31:0] _T_1154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1974;
  reg [31:0] _T_1154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1975;
  reg [31:0] _T_1155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1976;
  reg [31:0] _T_1155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1977;
  reg [31:0] _T_1156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1978;
  reg [31:0] _T_1156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1979;
  reg [31:0] _T_1157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1980;
  reg [31:0] _T_1157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1981;
  reg [31:0] _T_1158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1982;
  reg [31:0] _T_1158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1983;
  reg [31:0] _T_1159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1984;
  reg [31:0] _T_1159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1985;
  reg [31:0] _T_1160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1986;
  reg [31:0] _T_1160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1987;
  reg [31:0] _T_1161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1988;
  reg [31:0] _T_1161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1989;
  reg [31:0] _T_1162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1990;
  reg [31:0] _T_1162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1991;
  reg [31:0] _T_1163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1992;
  reg [31:0] _T_1163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1993;
  reg [31:0] _T_1164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1994;
  reg [31:0] _T_1164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1995;
  reg [31:0] _T_1165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1996;
  reg [31:0] _T_1165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1997;
  reg [31:0] _T_1166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1998;
  reg [31:0] _T_1166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1999;
  reg [31:0] _T_1167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2000;
  reg [31:0] _T_1167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2001;
  reg [31:0] _T_1168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2002;
  reg [31:0] _T_1168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2003;
  reg [31:0] _T_1169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2004;
  reg [31:0] _T_1169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2005;
  reg [31:0] _T_1170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2006;
  reg [31:0] _T_1170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2007;
  reg [31:0] _T_1171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2008;
  reg [31:0] _T_1171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2009;
  reg [31:0] _T_1172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2010;
  reg [31:0] _T_1172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2011;
  reg [31:0] _T_1173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2012;
  reg [31:0] _T_1173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2013;
  reg [31:0] _T_1174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2014;
  reg [31:0] _T_1174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2015;
  reg [31:0] _T_1175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2016;
  reg [31:0] _T_1175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2017;
  reg [31:0] _T_1176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2018;
  reg [31:0] _T_1176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2019;
  reg [31:0] _T_1177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2020;
  reg [31:0] _T_1177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2021;
  reg [31:0] _T_1178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2022;
  reg [31:0] _T_1178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2023;
  reg [31:0] _T_1179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2024;
  reg [31:0] _T_1179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2025;
  reg [31:0] _T_1180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2026;
  reg [31:0] _T_1180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2027;
  reg [31:0] _T_1181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2028;
  reg [31:0] _T_1181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2029;
  reg [31:0] _T_1182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2030;
  reg [31:0] _T_1182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2031;
  reg [31:0] _T_1183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2032;
  reg [31:0] _T_1183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2033;
  reg [31:0] _T_1184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2034;
  reg [31:0] _T_1184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2035;
  reg [31:0] _T_1185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2036;
  reg [31:0] _T_1185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2037;
  reg [31:0] _T_1186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2038;
  reg [31:0] _T_1186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2039;
  reg [31:0] _T_1187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2040;
  reg [31:0] _T_1187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2041;
  reg [31:0] _T_1188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2042;
  reg [31:0] _T_1188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2043;
  reg [31:0] _T_1189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2044;
  reg [31:0] _T_1189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2045;
  reg [31:0] _T_1190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2046;
  reg [31:0] _T_1190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2047;
  reg [31:0] _T_1191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2048;
  reg [31:0] _T_1191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2049;
  reg [31:0] _T_1194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2050;
  reg [31:0] _T_1194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2051;
  reg [31:0] _T_1195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2052;
  reg [31:0] _T_1195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2053;
  reg [31:0] _T_1196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2054;
  reg [31:0] _T_1196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2055;
  reg [31:0] _T_1197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2056;
  reg [31:0] _T_1197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2057;
  reg [31:0] _T_1198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2058;
  reg [31:0] _T_1198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2059;
  reg [31:0] _T_1199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2060;
  reg [31:0] _T_1199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2061;
  reg [31:0] _T_1200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2062;
  reg [31:0] _T_1200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2063;
  reg [31:0] _T_1201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2064;
  reg [31:0] _T_1201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2065;
  reg [31:0] _T_1202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2066;
  reg [31:0] _T_1202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2067;
  reg [31:0] _T_1203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2068;
  reg [31:0] _T_1203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2069;
  reg [31:0] _T_1204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2070;
  reg [31:0] _T_1204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2071;
  reg [31:0] _T_1205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2072;
  reg [31:0] _T_1205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2073;
  reg [31:0] _T_1206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2074;
  reg [31:0] _T_1206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2075;
  reg [31:0] _T_1207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2076;
  reg [31:0] _T_1207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2077;
  reg [31:0] _T_1208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2078;
  reg [31:0] _T_1208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2079;
  reg [31:0] _T_1209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2080;
  reg [31:0] _T_1209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2081;
  reg [31:0] _T_1210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2082;
  reg [31:0] _T_1210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2083;
  reg [31:0] _T_1211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2084;
  reg [31:0] _T_1211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2085;
  reg [31:0] _T_1212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2086;
  reg [31:0] _T_1212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2087;
  reg [31:0] _T_1213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2088;
  reg [31:0] _T_1213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2089;
  reg [31:0] _T_1214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2090;
  reg [31:0] _T_1214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2091;
  reg [31:0] _T_1215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2092;
  reg [31:0] _T_1215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2093;
  reg [31:0] _T_1216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2094;
  reg [31:0] _T_1216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2095;
  reg [31:0] _T_1217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2096;
  reg [31:0] _T_1217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2097;
  reg [31:0] _T_1218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2098;
  reg [31:0] _T_1218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2099;
  reg [31:0] _T_1219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2100;
  reg [31:0] _T_1219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2101;
  reg [31:0] _T_1220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2102;
  reg [31:0] _T_1220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2103;
  reg [31:0] _T_1221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2104;
  reg [31:0] _T_1221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2105;
  reg [31:0] _T_1222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2106;
  reg [31:0] _T_1222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2107;
  reg [31:0] _T_1223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2108;
  reg [31:0] _T_1223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2109;
  reg [31:0] _T_1224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2110;
  reg [31:0] _T_1224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2111;
  reg [31:0] _T_1225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2112;
  reg [31:0] _T_1225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2113;
  reg [31:0] _T_1226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2114;
  reg [31:0] _T_1226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2115;
  reg [31:0] _T_1227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2116;
  reg [31:0] _T_1227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2117;
  reg [31:0] _T_1228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2118;
  reg [31:0] _T_1228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2119;
  reg [31:0] _T_1229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2120;
  reg [31:0] _T_1229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2121;
  reg [31:0] _T_1230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2122;
  reg [31:0] _T_1230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2123;
  reg [31:0] _T_1231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2124;
  reg [31:0] _T_1231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2125;
  reg [31:0] _T_1232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2126;
  reg [31:0] _T_1232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2127;
  reg [31:0] _T_1233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2128;
  reg [31:0] _T_1233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2129;
  reg [31:0] _T_1234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2130;
  reg [31:0] _T_1234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2131;
  reg [31:0] _T_1235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2132;
  reg [31:0] _T_1235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2133;
  reg [31:0] _T_1236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2134;
  reg [31:0] _T_1236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2135;
  reg [31:0] _T_1237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2136;
  reg [31:0] _T_1237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2137;
  reg [31:0] _T_1238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2138;
  reg [31:0] _T_1238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2139;
  reg [31:0] _T_1239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2140;
  reg [31:0] _T_1239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2141;
  reg [31:0] _T_1240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2142;
  reg [31:0] _T_1240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2143;
  reg [31:0] _T_1241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2144;
  reg [31:0] _T_1241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2145;
  reg [31:0] _T_1242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2146;
  reg [31:0] _T_1242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2147;
  reg [31:0] _T_1243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2148;
  reg [31:0] _T_1243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2149;
  reg [31:0] _T_1244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2150;
  reg [31:0] _T_1244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2151;
  reg [31:0] _T_1245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2152;
  reg [31:0] _T_1245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2153;
  reg [31:0] _T_1246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2154;
  reg [31:0] _T_1246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2155;
  reg [31:0] _T_1247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2156;
  reg [31:0] _T_1247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2157;
  reg [31:0] _T_1248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2158;
  reg [31:0] _T_1248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2159;
  reg [31:0] _T_1249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2160;
  reg [31:0] _T_1249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2161;
  reg [31:0] _T_1250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2162;
  reg [31:0] _T_1250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2163;
  reg [31:0] _T_1251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2164;
  reg [31:0] _T_1251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2165;
  reg [31:0] _T_1252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2166;
  reg [31:0] _T_1252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2167;
  reg [31:0] _T_1253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2168;
  reg [31:0] _T_1253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2169;
  reg [31:0] _T_1254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2170;
  reg [31:0] _T_1254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2171;
  reg [31:0] _T_1255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2172;
  reg [31:0] _T_1255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2173;
  reg [31:0] _T_1256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2174;
  reg [31:0] _T_1256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2175;
  reg [31:0] _T_1257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2176;
  reg [31:0] _T_1257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2177;
  reg [31:0] _T_1258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2178;
  reg [31:0] _T_1258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2179;
  reg [31:0] _T_1259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2180;
  reg [31:0] _T_1259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2181;
  reg [31:0] _T_1260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2182;
  reg [31:0] _T_1260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2183;
  reg [31:0] _T_1261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2184;
  reg [31:0] _T_1261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2185;
  reg [31:0] _T_1262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2186;
  reg [31:0] _T_1262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2187;
  reg [31:0] _T_1263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2188;
  reg [31:0] _T_1263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2189;
  reg [31:0] _T_1264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2190;
  reg [31:0] _T_1264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2191;
  reg [31:0] _T_1265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2192;
  reg [31:0] _T_1265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2193;
  reg [31:0] _T_1266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2194;
  reg [31:0] _T_1266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2195;
  reg [31:0] _T_1267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2196;
  reg [31:0] _T_1267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2197;
  reg [31:0] _T_1268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2198;
  reg [31:0] _T_1268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2199;
  reg [31:0] _T_1269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2200;
  reg [31:0] _T_1269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2201;
  reg [31:0] _T_1270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2202;
  reg [31:0] _T_1270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2203;
  reg [31:0] _T_1271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2204;
  reg [31:0] _T_1271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2205;
  reg [31:0] _T_1272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2206;
  reg [31:0] _T_1272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2207;
  reg [31:0] _T_1273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2208;
  reg [31:0] _T_1273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2209;
  reg [31:0] _T_1274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2210;
  reg [31:0] _T_1274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2211;
  reg [31:0] _T_1275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2212;
  reg [31:0] _T_1275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2213;
  reg [31:0] _T_1276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2214;
  reg [31:0] _T_1276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2215;
  reg [31:0] _T_1277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2216;
  reg [31:0] _T_1277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2217;
  reg [31:0] _T_1278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2218;
  reg [31:0] _T_1278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2219;
  reg [31:0] _T_1279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2220;
  reg [31:0] _T_1279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2221;
  reg [31:0] _T_1280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2222;
  reg [31:0] _T_1280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2223;
  reg [31:0] _T_1281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2224;
  reg [31:0] _T_1281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2225;
  reg [31:0] _T_1282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2226;
  reg [31:0] _T_1282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2227;
  reg [31:0] _T_1283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2228;
  reg [31:0] _T_1283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2229;
  reg [31:0] _T_1284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2230;
  reg [31:0] _T_1284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2231;
  reg [31:0] _T_1285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2232;
  reg [31:0] _T_1285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2233;
  reg [31:0] _T_1286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2234;
  reg [31:0] _T_1286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2235;
  reg [31:0] _T_1287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2236;
  reg [31:0] _T_1287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2237;
  reg [31:0] _T_1288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2238;
  reg [31:0] _T_1288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2239;
  reg [31:0] _T_1289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2240;
  reg [31:0] _T_1289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2241;
  reg [31:0] _T_1290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2242;
  reg [31:0] _T_1290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2243;
  reg [31:0] _T_1291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2244;
  reg [31:0] _T_1291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2245;
  reg [31:0] _T_1292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2246;
  reg [31:0] _T_1292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2247;
  reg [31:0] _T_1293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2248;
  reg [31:0] _T_1293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2249;
  reg [31:0] _T_1294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2250;
  reg [31:0] _T_1294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2251;
  reg [31:0] _T_1295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2252;
  reg [31:0] _T_1295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2253;
  reg [31:0] _T_1296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2254;
  reg [31:0] _T_1296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2255;
  reg [31:0] _T_1297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2256;
  reg [31:0] _T_1297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2257;
  reg [31:0] _T_1298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2258;
  reg [31:0] _T_1298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2259;
  reg [31:0] _T_1299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2260;
  reg [31:0] _T_1299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2261;
  reg [31:0] _T_1300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2262;
  reg [31:0] _T_1300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2263;
  reg [31:0] _T_1301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2264;
  reg [31:0] _T_1301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2265;
  reg [31:0] _T_1302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2266;
  reg [31:0] _T_1302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2267;
  reg [31:0] _T_1303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2268;
  reg [31:0] _T_1303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2269;
  reg [31:0] _T_1304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2270;
  reg [31:0] _T_1304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2271;
  reg [31:0] _T_1305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2272;
  reg [31:0] _T_1305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2273;
  reg [31:0] _T_1306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2274;
  reg [31:0] _T_1306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2275;
  reg [31:0] _T_1307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2276;
  reg [31:0] _T_1307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2277;
  reg [31:0] _T_1308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2278;
  reg [31:0] _T_1308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2279;
  reg [31:0] _T_1309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2280;
  reg [31:0] _T_1309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2281;
  reg [31:0] _T_1310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2282;
  reg [31:0] _T_1310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2283;
  reg [31:0] _T_1311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2284;
  reg [31:0] _T_1311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2285;
  reg [31:0] _T_1312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2286;
  reg [31:0] _T_1312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2287;
  reg [31:0] _T_1313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2288;
  reg [31:0] _T_1313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2289;
  reg [31:0] _T_1314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2290;
  reg [31:0] _T_1314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2291;
  reg [31:0] _T_1315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2292;
  reg [31:0] _T_1315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2293;
  reg [31:0] _T_1316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2294;
  reg [31:0] _T_1316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2295;
  reg [31:0] _T_1317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2296;
  reg [31:0] _T_1317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2297;
  reg [31:0] _T_1318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2298;
  reg [31:0] _T_1318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2299;
  reg [31:0] _T_1319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2300;
  reg [31:0] _T_1319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2301;
  reg [31:0] _T_1320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2302;
  reg [31:0] _T_1320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2303;
  reg [31:0] _T_1321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2304;
  reg [31:0] _T_1321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2305;
  wire [31:0] _GEN_3842; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3843; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3844; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3845; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3846; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3847; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3848; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3849; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3850; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3851; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3852; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3853; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3854; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3855; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3856; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3857; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3858; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3859; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3860; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3861; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3862; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3863; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3864; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3865; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3866; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3867; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3868; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3869; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3870; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3871; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3872; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3873; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3874; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3875; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3876; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3877; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3878; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3879; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3880; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3881; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3882; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3883; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3884; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3885; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3886; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3887; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3888; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3889; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3890; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3891; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3892; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3893; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3894; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3895; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3896; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3897; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3898; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3899; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3900; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3901; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3902; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3903; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3904; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3905; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3906; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3907; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3908; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3909; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3910; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3911; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3912; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3913; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3914; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3915; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3916; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3917; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3918; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3919; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3920; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3921; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3922; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3923; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3924; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3925; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3926; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3927; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3928; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3929; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3930; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3931; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3932; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3933; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3934; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3935; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3936; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3937; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3938; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3939; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3940; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3941; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3942; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3943; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3944; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3945; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3946; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3947; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3948; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3949; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3950; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3951; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3952; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3953; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3954; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3955; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3956; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3957; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3958; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3959; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3960; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3961; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3962; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3963; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3964; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3965; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3966; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3967; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3970; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3971; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3972; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3973; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3974; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3975; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3976; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3977; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3978; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3979; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3980; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3981; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3982; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3983; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3984; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3985; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3986; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3987; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3988; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3989; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3990; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3991; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3992; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3993; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3994; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3995; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3996; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3997; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3998; // @[FFT.scala 35:12]
  wire [31:0] _GEN_3999; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4000; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4001; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4002; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4003; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4004; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4005; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4006; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4007; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4008; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4009; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4010; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4011; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4012; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4013; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4014; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4015; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4016; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4017; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4018; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4019; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4020; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4021; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4022; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4023; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4024; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4025; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4026; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4027; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4028; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4029; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4030; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4031; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4032; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4033; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4034; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4035; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4036; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4037; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4038; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4039; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4040; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4041; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4042; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4043; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4044; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4045; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4046; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4047; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4048; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4049; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4050; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4051; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4052; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4053; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4054; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4055; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4056; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4057; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4058; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4059; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4060; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4061; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4062; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4063; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4064; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4065; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4066; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4067; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4068; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4069; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4070; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4071; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4072; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4073; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4074; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4075; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4076; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4077; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4078; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4079; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4080; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4081; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4082; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4083; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4084; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4085; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4086; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4087; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4088; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4089; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4090; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4091; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4092; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4093; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4094; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4095; // @[FFT.scala 35:12]
  reg [31:0] _T_1327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2306;
  reg [31:0] _T_1327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2307;
  reg [31:0] _T_1328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2308;
  reg [31:0] _T_1328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2309;
  reg [31:0] _T_1329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2310;
  reg [31:0] _T_1329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2311;
  reg [31:0] _T_1330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2312;
  reg [31:0] _T_1330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2313;
  reg [31:0] _T_1331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2314;
  reg [31:0] _T_1331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2315;
  reg [31:0] _T_1332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2316;
  reg [31:0] _T_1332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2317;
  reg [31:0] _T_1333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2318;
  reg [31:0] _T_1333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2319;
  reg [31:0] _T_1334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2320;
  reg [31:0] _T_1334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2321;
  reg [31:0] _T_1335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2322;
  reg [31:0] _T_1335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2323;
  reg [31:0] _T_1336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2324;
  reg [31:0] _T_1336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2325;
  reg [31:0] _T_1337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2326;
  reg [31:0] _T_1337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2327;
  reg [31:0] _T_1338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2328;
  reg [31:0] _T_1338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2329;
  reg [31:0] _T_1339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2330;
  reg [31:0] _T_1339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2331;
  reg [31:0] _T_1340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2332;
  reg [31:0] _T_1340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2333;
  reg [31:0] _T_1341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2334;
  reg [31:0] _T_1341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2335;
  reg [31:0] _T_1342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2336;
  reg [31:0] _T_1342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2337;
  reg [31:0] _T_1343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2338;
  reg [31:0] _T_1343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2339;
  reg [31:0] _T_1344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2340;
  reg [31:0] _T_1344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2341;
  reg [31:0] _T_1345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2342;
  reg [31:0] _T_1345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2343;
  reg [31:0] _T_1346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2344;
  reg [31:0] _T_1346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2345;
  reg [31:0] _T_1347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2346;
  reg [31:0] _T_1347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2347;
  reg [31:0] _T_1348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2348;
  reg [31:0] _T_1348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2349;
  reg [31:0] _T_1349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2350;
  reg [31:0] _T_1349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2351;
  reg [31:0] _T_1350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2352;
  reg [31:0] _T_1350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2353;
  reg [31:0] _T_1351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2354;
  reg [31:0] _T_1351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2355;
  reg [31:0] _T_1352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2356;
  reg [31:0] _T_1352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2357;
  reg [31:0] _T_1353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2358;
  reg [31:0] _T_1353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2359;
  reg [31:0] _T_1354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2360;
  reg [31:0] _T_1354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2361;
  reg [31:0] _T_1355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2362;
  reg [31:0] _T_1355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2363;
  reg [31:0] _T_1356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2364;
  reg [31:0] _T_1356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2365;
  reg [31:0] _T_1357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2366;
  reg [31:0] _T_1357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2367;
  reg [31:0] _T_1358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2368;
  reg [31:0] _T_1358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2369;
  reg [31:0] _T_1359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2370;
  reg [31:0] _T_1359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2371;
  reg [31:0] _T_1360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2372;
  reg [31:0] _T_1360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2373;
  reg [31:0] _T_1361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2374;
  reg [31:0] _T_1361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2375;
  reg [31:0] _T_1362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2376;
  reg [31:0] _T_1362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2377;
  reg [31:0] _T_1363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2378;
  reg [31:0] _T_1363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2379;
  reg [31:0] _T_1364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2380;
  reg [31:0] _T_1364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2381;
  reg [31:0] _T_1365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2382;
  reg [31:0] _T_1365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2383;
  reg [31:0] _T_1366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2384;
  reg [31:0] _T_1366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2385;
  reg [31:0] _T_1367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2386;
  reg [31:0] _T_1367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2387;
  reg [31:0] _T_1368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2388;
  reg [31:0] _T_1368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2389;
  reg [31:0] _T_1369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2390;
  reg [31:0] _T_1369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2391;
  reg [31:0] _T_1370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2392;
  reg [31:0] _T_1370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2393;
  reg [31:0] _T_1371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2394;
  reg [31:0] _T_1371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2395;
  reg [31:0] _T_1372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2396;
  reg [31:0] _T_1372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2397;
  reg [31:0] _T_1373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2398;
  reg [31:0] _T_1373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2399;
  reg [31:0] _T_1374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2400;
  reg [31:0] _T_1374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2401;
  reg [31:0] _T_1375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2402;
  reg [31:0] _T_1375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2403;
  reg [31:0] _T_1376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2404;
  reg [31:0] _T_1376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2405;
  reg [31:0] _T_1377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2406;
  reg [31:0] _T_1377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2407;
  reg [31:0] _T_1378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2408;
  reg [31:0] _T_1378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2409;
  reg [31:0] _T_1379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2410;
  reg [31:0] _T_1379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2411;
  reg [31:0] _T_1380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2412;
  reg [31:0] _T_1380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2413;
  reg [31:0] _T_1381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2414;
  reg [31:0] _T_1381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2415;
  reg [31:0] _T_1382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2416;
  reg [31:0] _T_1382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2417;
  reg [31:0] _T_1383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2418;
  reg [31:0] _T_1383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2419;
  reg [31:0] _T_1384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2420;
  reg [31:0] _T_1384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2421;
  reg [31:0] _T_1385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2422;
  reg [31:0] _T_1385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2423;
  reg [31:0] _T_1386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2424;
  reg [31:0] _T_1386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2425;
  reg [31:0] _T_1387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2426;
  reg [31:0] _T_1387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2427;
  reg [31:0] _T_1388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2428;
  reg [31:0] _T_1388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2429;
  reg [31:0] _T_1389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2430;
  reg [31:0] _T_1389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2431;
  reg [31:0] _T_1390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2432;
  reg [31:0] _T_1390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2433;
  reg [31:0] _T_1391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2434;
  reg [31:0] _T_1391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2435;
  reg [31:0] _T_1392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2436;
  reg [31:0] _T_1392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2437;
  reg [31:0] _T_1393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2438;
  reg [31:0] _T_1393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2439;
  reg [31:0] _T_1394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2440;
  reg [31:0] _T_1394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2441;
  reg [31:0] _T_1395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2442;
  reg [31:0] _T_1395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2443;
  reg [31:0] _T_1396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2444;
  reg [31:0] _T_1396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2445;
  reg [31:0] _T_1397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2446;
  reg [31:0] _T_1397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2447;
  reg [31:0] _T_1398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2448;
  reg [31:0] _T_1398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2449;
  reg [31:0] _T_1399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2450;
  reg [31:0] _T_1399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2451;
  reg [31:0] _T_1400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2452;
  reg [31:0] _T_1400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2453;
  reg [31:0] _T_1401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2454;
  reg [31:0] _T_1401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2455;
  reg [31:0] _T_1402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2456;
  reg [31:0] _T_1402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2457;
  reg [31:0] _T_1403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2458;
  reg [31:0] _T_1403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2459;
  reg [31:0] _T_1404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2460;
  reg [31:0] _T_1404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2461;
  reg [31:0] _T_1405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2462;
  reg [31:0] _T_1405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2463;
  reg [31:0] _T_1406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2464;
  reg [31:0] _T_1406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2465;
  reg [31:0] _T_1407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2466;
  reg [31:0] _T_1407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2467;
  reg [31:0] _T_1408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2468;
  reg [31:0] _T_1408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2469;
  reg [31:0] _T_1409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2470;
  reg [31:0] _T_1409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2471;
  reg [31:0] _T_1410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2472;
  reg [31:0] _T_1410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2473;
  reg [31:0] _T_1411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2474;
  reg [31:0] _T_1411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2475;
  reg [31:0] _T_1412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2476;
  reg [31:0] _T_1412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2477;
  reg [31:0] _T_1413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2478;
  reg [31:0] _T_1413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2479;
  reg [31:0] _T_1414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2480;
  reg [31:0] _T_1414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2481;
  reg [31:0] _T_1415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2482;
  reg [31:0] _T_1415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2483;
  reg [31:0] _T_1416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2484;
  reg [31:0] _T_1416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2485;
  reg [31:0] _T_1417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2486;
  reg [31:0] _T_1417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2487;
  reg [31:0] _T_1418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2488;
  reg [31:0] _T_1418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2489;
  reg [31:0] _T_1419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2490;
  reg [31:0] _T_1419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2491;
  reg [31:0] _T_1420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2492;
  reg [31:0] _T_1420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2493;
  reg [31:0] _T_1421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2494;
  reg [31:0] _T_1421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2495;
  reg [31:0] _T_1422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2496;
  reg [31:0] _T_1422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2497;
  reg [31:0] _T_1423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2498;
  reg [31:0] _T_1423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2499;
  reg [31:0] _T_1424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2500;
  reg [31:0] _T_1424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2501;
  reg [31:0] _T_1425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2502;
  reg [31:0] _T_1425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2503;
  reg [31:0] _T_1426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2504;
  reg [31:0] _T_1426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2505;
  reg [31:0] _T_1427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2506;
  reg [31:0] _T_1427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2507;
  reg [31:0] _T_1428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2508;
  reg [31:0] _T_1428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2509;
  reg [31:0] _T_1429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2510;
  reg [31:0] _T_1429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2511;
  reg [31:0] _T_1430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2512;
  reg [31:0] _T_1430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2513;
  reg [31:0] _T_1431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2514;
  reg [31:0] _T_1431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2515;
  reg [31:0] _T_1432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2516;
  reg [31:0] _T_1432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2517;
  reg [31:0] _T_1433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2518;
  reg [31:0] _T_1433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2519;
  reg [31:0] _T_1434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2520;
  reg [31:0] _T_1434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2521;
  reg [31:0] _T_1435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2522;
  reg [31:0] _T_1435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2523;
  reg [31:0] _T_1436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2524;
  reg [31:0] _T_1436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2525;
  reg [31:0] _T_1437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2526;
  reg [31:0] _T_1437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2527;
  reg [31:0] _T_1438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2528;
  reg [31:0] _T_1438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2529;
  reg [31:0] _T_1439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2530;
  reg [31:0] _T_1439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2531;
  reg [31:0] _T_1440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2532;
  reg [31:0] _T_1440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2533;
  reg [31:0] _T_1441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2534;
  reg [31:0] _T_1441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2535;
  reg [31:0] _T_1442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2536;
  reg [31:0] _T_1442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2537;
  reg [31:0] _T_1443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2538;
  reg [31:0] _T_1443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2539;
  reg [31:0] _T_1444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2540;
  reg [31:0] _T_1444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2541;
  reg [31:0] _T_1445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2542;
  reg [31:0] _T_1445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2543;
  reg [31:0] _T_1446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2544;
  reg [31:0] _T_1446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2545;
  reg [31:0] _T_1447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2546;
  reg [31:0] _T_1447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2547;
  reg [31:0] _T_1448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2548;
  reg [31:0] _T_1448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2549;
  reg [31:0] _T_1449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2550;
  reg [31:0] _T_1449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2551;
  reg [31:0] _T_1450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2552;
  reg [31:0] _T_1450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2553;
  reg [31:0] _T_1451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2554;
  reg [31:0] _T_1451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2555;
  reg [31:0] _T_1452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2556;
  reg [31:0] _T_1452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2557;
  reg [31:0] _T_1453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2558;
  reg [31:0] _T_1453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2559;
  reg [31:0] _T_1454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2560;
  reg [31:0] _T_1454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2561;
  reg [31:0] _T_1457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2562;
  reg [31:0] _T_1457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2563;
  reg [31:0] _T_1458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2564;
  reg [31:0] _T_1458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2565;
  reg [31:0] _T_1459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2566;
  reg [31:0] _T_1459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2567;
  reg [31:0] _T_1460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2568;
  reg [31:0] _T_1460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2569;
  reg [31:0] _T_1461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2570;
  reg [31:0] _T_1461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2571;
  reg [31:0] _T_1462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2572;
  reg [31:0] _T_1462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2573;
  reg [31:0] _T_1463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2574;
  reg [31:0] _T_1463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2575;
  reg [31:0] _T_1464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2576;
  reg [31:0] _T_1464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2577;
  reg [31:0] _T_1465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2578;
  reg [31:0] _T_1465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2579;
  reg [31:0] _T_1466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2580;
  reg [31:0] _T_1466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2581;
  reg [31:0] _T_1467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2582;
  reg [31:0] _T_1467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2583;
  reg [31:0] _T_1468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2584;
  reg [31:0] _T_1468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2585;
  reg [31:0] _T_1469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2586;
  reg [31:0] _T_1469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2587;
  reg [31:0] _T_1470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2588;
  reg [31:0] _T_1470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2589;
  reg [31:0] _T_1471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2590;
  reg [31:0] _T_1471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2591;
  reg [31:0] _T_1472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2592;
  reg [31:0] _T_1472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2593;
  reg [31:0] _T_1473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2594;
  reg [31:0] _T_1473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2595;
  reg [31:0] _T_1474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2596;
  reg [31:0] _T_1474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2597;
  reg [31:0] _T_1475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2598;
  reg [31:0] _T_1475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2599;
  reg [31:0] _T_1476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2600;
  reg [31:0] _T_1476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2601;
  reg [31:0] _T_1477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2602;
  reg [31:0] _T_1477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2603;
  reg [31:0] _T_1478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2604;
  reg [31:0] _T_1478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2605;
  reg [31:0] _T_1479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2606;
  reg [31:0] _T_1479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2607;
  reg [31:0] _T_1480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2608;
  reg [31:0] _T_1480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2609;
  reg [31:0] _T_1481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2610;
  reg [31:0] _T_1481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2611;
  reg [31:0] _T_1482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2612;
  reg [31:0] _T_1482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2613;
  reg [31:0] _T_1483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2614;
  reg [31:0] _T_1483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2615;
  reg [31:0] _T_1484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2616;
  reg [31:0] _T_1484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2617;
  reg [31:0] _T_1485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2618;
  reg [31:0] _T_1485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2619;
  reg [31:0] _T_1486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2620;
  reg [31:0] _T_1486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2621;
  reg [31:0] _T_1487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2622;
  reg [31:0] _T_1487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2623;
  reg [31:0] _T_1488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2624;
  reg [31:0] _T_1488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2625;
  reg [31:0] _T_1489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2626;
  reg [31:0] _T_1489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2627;
  reg [31:0] _T_1490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2628;
  reg [31:0] _T_1490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2629;
  reg [31:0] _T_1491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2630;
  reg [31:0] _T_1491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2631;
  reg [31:0] _T_1492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2632;
  reg [31:0] _T_1492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2633;
  reg [31:0] _T_1493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2634;
  reg [31:0] _T_1493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2635;
  reg [31:0] _T_1494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2636;
  reg [31:0] _T_1494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2637;
  reg [31:0] _T_1495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2638;
  reg [31:0] _T_1495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2639;
  reg [31:0] _T_1496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2640;
  reg [31:0] _T_1496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2641;
  reg [31:0] _T_1497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2642;
  reg [31:0] _T_1497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2643;
  reg [31:0] _T_1498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2644;
  reg [31:0] _T_1498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2645;
  reg [31:0] _T_1499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2646;
  reg [31:0] _T_1499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2647;
  reg [31:0] _T_1500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2648;
  reg [31:0] _T_1500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2649;
  reg [31:0] _T_1501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2650;
  reg [31:0] _T_1501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2651;
  reg [31:0] _T_1502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2652;
  reg [31:0] _T_1502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2653;
  reg [31:0] _T_1503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2654;
  reg [31:0] _T_1503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2655;
  reg [31:0] _T_1504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2656;
  reg [31:0] _T_1504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2657;
  reg [31:0] _T_1505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2658;
  reg [31:0] _T_1505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2659;
  reg [31:0] _T_1506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2660;
  reg [31:0] _T_1506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2661;
  reg [31:0] _T_1507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2662;
  reg [31:0] _T_1507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2663;
  reg [31:0] _T_1508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2664;
  reg [31:0] _T_1508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2665;
  reg [31:0] _T_1509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2666;
  reg [31:0] _T_1509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2667;
  reg [31:0] _T_1510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2668;
  reg [31:0] _T_1510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2669;
  reg [31:0] _T_1511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2670;
  reg [31:0] _T_1511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2671;
  reg [31:0] _T_1512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2672;
  reg [31:0] _T_1512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2673;
  reg [31:0] _T_1513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2674;
  reg [31:0] _T_1513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2675;
  reg [31:0] _T_1514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2676;
  reg [31:0] _T_1514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2677;
  reg [31:0] _T_1515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2678;
  reg [31:0] _T_1515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2679;
  reg [31:0] _T_1516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2680;
  reg [31:0] _T_1516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2681;
  reg [31:0] _T_1517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2682;
  reg [31:0] _T_1517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2683;
  reg [31:0] _T_1518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2684;
  reg [31:0] _T_1518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2685;
  reg [31:0] _T_1519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2686;
  reg [31:0] _T_1519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2687;
  reg [31:0] _T_1520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2688;
  reg [31:0] _T_1520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2689;
  wire [31:0] _GEN_4482; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4483; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4484; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4485; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4486; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4487; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4488; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4489; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4490; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4491; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4492; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4493; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4494; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4495; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4496; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4497; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4498; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4499; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4500; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4501; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4502; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4503; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4504; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4505; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4506; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4507; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4508; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4509; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4510; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4511; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4512; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4513; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4514; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4515; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4516; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4517; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4518; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4519; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4520; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4521; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4522; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4523; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4524; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4525; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4526; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4527; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4528; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4529; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4530; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4531; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4532; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4533; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4534; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4535; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4536; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4537; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4538; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4539; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4540; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4541; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4542; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4543; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4546; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4547; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4548; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4549; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4550; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4551; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4552; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4553; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4554; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4555; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4556; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4557; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4558; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4559; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4560; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4561; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4562; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4563; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4564; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4565; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4566; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4567; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4568; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4569; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4570; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4571; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4572; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4573; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4574; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4575; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4576; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4577; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4578; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4579; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4580; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4581; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4582; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4583; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4584; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4585; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4586; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4587; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4588; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4589; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4590; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4591; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4592; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4593; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4594; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4595; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4596; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4597; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4598; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4599; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4600; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4601; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4602; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4603; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4604; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4605; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4606; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4607; // @[FFT.scala 35:12]
  reg [31:0] _T_1526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2690;
  reg [31:0] _T_1526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2691;
  reg [31:0] _T_1527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2692;
  reg [31:0] _T_1527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2693;
  reg [31:0] _T_1528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2694;
  reg [31:0] _T_1528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2695;
  reg [31:0] _T_1529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2696;
  reg [31:0] _T_1529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2697;
  reg [31:0] _T_1530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2698;
  reg [31:0] _T_1530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2699;
  reg [31:0] _T_1531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2700;
  reg [31:0] _T_1531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2701;
  reg [31:0] _T_1532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2702;
  reg [31:0] _T_1532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2703;
  reg [31:0] _T_1533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2704;
  reg [31:0] _T_1533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2705;
  reg [31:0] _T_1534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2706;
  reg [31:0] _T_1534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2707;
  reg [31:0] _T_1535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2708;
  reg [31:0] _T_1535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2709;
  reg [31:0] _T_1536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2710;
  reg [31:0] _T_1536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2711;
  reg [31:0] _T_1537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2712;
  reg [31:0] _T_1537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2713;
  reg [31:0] _T_1538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2714;
  reg [31:0] _T_1538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2715;
  reg [31:0] _T_1539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2716;
  reg [31:0] _T_1539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2717;
  reg [31:0] _T_1540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2718;
  reg [31:0] _T_1540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2719;
  reg [31:0] _T_1541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2720;
  reg [31:0] _T_1541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2721;
  reg [31:0] _T_1542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2722;
  reg [31:0] _T_1542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2723;
  reg [31:0] _T_1543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2724;
  reg [31:0] _T_1543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2725;
  reg [31:0] _T_1544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2726;
  reg [31:0] _T_1544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2727;
  reg [31:0] _T_1545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2728;
  reg [31:0] _T_1545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2729;
  reg [31:0] _T_1546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2730;
  reg [31:0] _T_1546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2731;
  reg [31:0] _T_1547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2732;
  reg [31:0] _T_1547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2733;
  reg [31:0] _T_1548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2734;
  reg [31:0] _T_1548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2735;
  reg [31:0] _T_1549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2736;
  reg [31:0] _T_1549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2737;
  reg [31:0] _T_1550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2738;
  reg [31:0] _T_1550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2739;
  reg [31:0] _T_1551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2740;
  reg [31:0] _T_1551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2741;
  reg [31:0] _T_1552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2742;
  reg [31:0] _T_1552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2743;
  reg [31:0] _T_1553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2744;
  reg [31:0] _T_1553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2745;
  reg [31:0] _T_1554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2746;
  reg [31:0] _T_1554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2747;
  reg [31:0] _T_1555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2748;
  reg [31:0] _T_1555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2749;
  reg [31:0] _T_1556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2750;
  reg [31:0] _T_1556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2751;
  reg [31:0] _T_1557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2752;
  reg [31:0] _T_1557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2753;
  reg [31:0] _T_1558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2754;
  reg [31:0] _T_1558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2755;
  reg [31:0] _T_1559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2756;
  reg [31:0] _T_1559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2757;
  reg [31:0] _T_1560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2758;
  reg [31:0] _T_1560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2759;
  reg [31:0] _T_1561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2760;
  reg [31:0] _T_1561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2761;
  reg [31:0] _T_1562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2762;
  reg [31:0] _T_1562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2763;
  reg [31:0] _T_1563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2764;
  reg [31:0] _T_1563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2765;
  reg [31:0] _T_1564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2766;
  reg [31:0] _T_1564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2767;
  reg [31:0] _T_1565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2768;
  reg [31:0] _T_1565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2769;
  reg [31:0] _T_1566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2770;
  reg [31:0] _T_1566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2771;
  reg [31:0] _T_1567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2772;
  reg [31:0] _T_1567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2773;
  reg [31:0] _T_1568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2774;
  reg [31:0] _T_1568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2775;
  reg [31:0] _T_1569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2776;
  reg [31:0] _T_1569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2777;
  reg [31:0] _T_1570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2778;
  reg [31:0] _T_1570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2779;
  reg [31:0] _T_1571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2780;
  reg [31:0] _T_1571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2781;
  reg [31:0] _T_1572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2782;
  reg [31:0] _T_1572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2783;
  reg [31:0] _T_1573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2784;
  reg [31:0] _T_1573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2785;
  reg [31:0] _T_1574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2786;
  reg [31:0] _T_1574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2787;
  reg [31:0] _T_1575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2788;
  reg [31:0] _T_1575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2789;
  reg [31:0] _T_1576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2790;
  reg [31:0] _T_1576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2791;
  reg [31:0] _T_1577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2792;
  reg [31:0] _T_1577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2793;
  reg [31:0] _T_1578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2794;
  reg [31:0] _T_1578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2795;
  reg [31:0] _T_1579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2796;
  reg [31:0] _T_1579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2797;
  reg [31:0] _T_1580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2798;
  reg [31:0] _T_1580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2799;
  reg [31:0] _T_1581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2800;
  reg [31:0] _T_1581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2801;
  reg [31:0] _T_1582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2802;
  reg [31:0] _T_1582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2803;
  reg [31:0] _T_1583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2804;
  reg [31:0] _T_1583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2805;
  reg [31:0] _T_1584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2806;
  reg [31:0] _T_1584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2807;
  reg [31:0] _T_1585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2808;
  reg [31:0] _T_1585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2809;
  reg [31:0] _T_1586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2810;
  reg [31:0] _T_1586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2811;
  reg [31:0] _T_1587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2812;
  reg [31:0] _T_1587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2813;
  reg [31:0] _T_1588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2814;
  reg [31:0] _T_1588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2815;
  reg [31:0] _T_1589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2816;
  reg [31:0] _T_1589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2817;
  reg [31:0] _T_1592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2818;
  reg [31:0] _T_1592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2819;
  reg [31:0] _T_1593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2820;
  reg [31:0] _T_1593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2821;
  reg [31:0] _T_1594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2822;
  reg [31:0] _T_1594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2823;
  reg [31:0] _T_1595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2824;
  reg [31:0] _T_1595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2825;
  reg [31:0] _T_1596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2826;
  reg [31:0] _T_1596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2827;
  reg [31:0] _T_1597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2828;
  reg [31:0] _T_1597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2829;
  reg [31:0] _T_1598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2830;
  reg [31:0] _T_1598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2831;
  reg [31:0] _T_1599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2832;
  reg [31:0] _T_1599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2833;
  reg [31:0] _T_1600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2834;
  reg [31:0] _T_1600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2835;
  reg [31:0] _T_1601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2836;
  reg [31:0] _T_1601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2837;
  reg [31:0] _T_1602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2838;
  reg [31:0] _T_1602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2839;
  reg [31:0] _T_1603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2840;
  reg [31:0] _T_1603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2841;
  reg [31:0] _T_1604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2842;
  reg [31:0] _T_1604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2843;
  reg [31:0] _T_1605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2844;
  reg [31:0] _T_1605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2845;
  reg [31:0] _T_1606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2846;
  reg [31:0] _T_1606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2847;
  reg [31:0] _T_1607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2848;
  reg [31:0] _T_1607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2849;
  reg [31:0] _T_1608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2850;
  reg [31:0] _T_1608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2851;
  reg [31:0] _T_1609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2852;
  reg [31:0] _T_1609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2853;
  reg [31:0] _T_1610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2854;
  reg [31:0] _T_1610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2855;
  reg [31:0] _T_1611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2856;
  reg [31:0] _T_1611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2857;
  reg [31:0] _T_1612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2858;
  reg [31:0] _T_1612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2859;
  reg [31:0] _T_1613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2860;
  reg [31:0] _T_1613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2861;
  reg [31:0] _T_1614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2862;
  reg [31:0] _T_1614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2863;
  reg [31:0] _T_1615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2864;
  reg [31:0] _T_1615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2865;
  reg [31:0] _T_1616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2866;
  reg [31:0] _T_1616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2867;
  reg [31:0] _T_1617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2868;
  reg [31:0] _T_1617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2869;
  reg [31:0] _T_1618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2870;
  reg [31:0] _T_1618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2871;
  reg [31:0] _T_1619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2872;
  reg [31:0] _T_1619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2873;
  reg [31:0] _T_1620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2874;
  reg [31:0] _T_1620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2875;
  reg [31:0] _T_1621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2876;
  reg [31:0] _T_1621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2877;
  reg [31:0] _T_1622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2878;
  reg [31:0] _T_1622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2879;
  reg [31:0] _T_1623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2880;
  reg [31:0] _T_1623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2881;
  wire [31:0] _GEN_4802; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4803; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4804; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4805; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4806; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4807; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4808; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4809; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4810; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4811; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4812; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4813; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4814; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4815; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4816; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4817; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4818; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4819; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4820; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4821; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4822; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4823; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4824; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4825; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4826; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4827; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4828; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4829; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4830; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4831; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4834; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4835; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4836; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4837; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4838; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4839; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4840; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4841; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4842; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4843; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4844; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4845; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4846; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4847; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4848; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4849; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4850; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4851; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4852; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4853; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4854; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4855; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4856; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4857; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4858; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4859; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4860; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4861; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4862; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4863; // @[FFT.scala 35:12]
  reg [31:0] _T_1629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2882;
  reg [31:0] _T_1629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2883;
  reg [31:0] _T_1630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2884;
  reg [31:0] _T_1630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2885;
  reg [31:0] _T_1631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2886;
  reg [31:0] _T_1631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2887;
  reg [31:0] _T_1632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2888;
  reg [31:0] _T_1632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2889;
  reg [31:0] _T_1633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2890;
  reg [31:0] _T_1633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2891;
  reg [31:0] _T_1634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2892;
  reg [31:0] _T_1634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2893;
  reg [31:0] _T_1635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2894;
  reg [31:0] _T_1635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2895;
  reg [31:0] _T_1636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2896;
  reg [31:0] _T_1636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2897;
  reg [31:0] _T_1637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2898;
  reg [31:0] _T_1637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2899;
  reg [31:0] _T_1638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2900;
  reg [31:0] _T_1638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2901;
  reg [31:0] _T_1639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2902;
  reg [31:0] _T_1639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2903;
  reg [31:0] _T_1640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2904;
  reg [31:0] _T_1640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2905;
  reg [31:0] _T_1641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2906;
  reg [31:0] _T_1641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2907;
  reg [31:0] _T_1642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2908;
  reg [31:0] _T_1642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2909;
  reg [31:0] _T_1643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2910;
  reg [31:0] _T_1643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2911;
  reg [31:0] _T_1644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2912;
  reg [31:0] _T_1644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2913;
  reg [31:0] _T_1645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2914;
  reg [31:0] _T_1645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2915;
  reg [31:0] _T_1646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2916;
  reg [31:0] _T_1646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2917;
  reg [31:0] _T_1647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2918;
  reg [31:0] _T_1647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2919;
  reg [31:0] _T_1648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2920;
  reg [31:0] _T_1648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2921;
  reg [31:0] _T_1649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2922;
  reg [31:0] _T_1649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2923;
  reg [31:0] _T_1650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2924;
  reg [31:0] _T_1650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2925;
  reg [31:0] _T_1651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2926;
  reg [31:0] _T_1651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2927;
  reg [31:0] _T_1652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2928;
  reg [31:0] _T_1652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2929;
  reg [31:0] _T_1653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2930;
  reg [31:0] _T_1653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2931;
  reg [31:0] _T_1654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2932;
  reg [31:0] _T_1654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2933;
  reg [31:0] _T_1655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2934;
  reg [31:0] _T_1655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2935;
  reg [31:0] _T_1656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2936;
  reg [31:0] _T_1656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2937;
  reg [31:0] _T_1657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2938;
  reg [31:0] _T_1657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2939;
  reg [31:0] _T_1658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2940;
  reg [31:0] _T_1658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2941;
  reg [31:0] _T_1659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2942;
  reg [31:0] _T_1659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2943;
  reg [31:0] _T_1660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2944;
  reg [31:0] _T_1660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2945;
  reg [31:0] _T_1663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2946;
  reg [31:0] _T_1663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2947;
  reg [31:0] _T_1664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2948;
  reg [31:0] _T_1664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2949;
  reg [31:0] _T_1665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2950;
  reg [31:0] _T_1665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2951;
  reg [31:0] _T_1666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2952;
  reg [31:0] _T_1666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2953;
  reg [31:0] _T_1667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2954;
  reg [31:0] _T_1667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2955;
  reg [31:0] _T_1668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2956;
  reg [31:0] _T_1668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2957;
  reg [31:0] _T_1669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2958;
  reg [31:0] _T_1669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2959;
  reg [31:0] _T_1670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2960;
  reg [31:0] _T_1670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2961;
  reg [31:0] _T_1671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2962;
  reg [31:0] _T_1671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2963;
  reg [31:0] _T_1672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2964;
  reg [31:0] _T_1672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2965;
  reg [31:0] _T_1673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2966;
  reg [31:0] _T_1673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2967;
  reg [31:0] _T_1674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2968;
  reg [31:0] _T_1674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2969;
  reg [31:0] _T_1675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2970;
  reg [31:0] _T_1675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2971;
  reg [31:0] _T_1676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2972;
  reg [31:0] _T_1676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2973;
  reg [31:0] _T_1677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2974;
  reg [31:0] _T_1677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2975;
  reg [31:0] _T_1678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2976;
  reg [31:0] _T_1678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2977;
  wire [31:0] _GEN_4962; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4963; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4964; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4965; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4966; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4967; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4968; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4969; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4970; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4971; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4972; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4973; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4974; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4975; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4978; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4979; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4980; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4981; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4982; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4983; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4984; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4985; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4986; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4987; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4988; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4989; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4990; // @[FFT.scala 35:12]
  wire [31:0] _GEN_4991; // @[FFT.scala 35:12]
  reg [31:0] _T_1684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2978;
  reg [31:0] _T_1684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2979;
  reg [31:0] _T_1685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2980;
  reg [31:0] _T_1685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2981;
  reg [31:0] _T_1686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2982;
  reg [31:0] _T_1686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2983;
  reg [31:0] _T_1687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2984;
  reg [31:0] _T_1687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2985;
  reg [31:0] _T_1688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2986;
  reg [31:0] _T_1688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2987;
  reg [31:0] _T_1689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2988;
  reg [31:0] _T_1689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2989;
  reg [31:0] _T_1690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2990;
  reg [31:0] _T_1690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2991;
  reg [31:0] _T_1691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2992;
  reg [31:0] _T_1691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2993;
  reg [31:0] _T_1692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2994;
  reg [31:0] _T_1692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2995;
  reg [31:0] _T_1693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2996;
  reg [31:0] _T_1693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2997;
  reg [31:0] _T_1694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2998;
  reg [31:0] _T_1694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2999;
  reg [31:0] _T_1695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3000;
  reg [31:0] _T_1695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3001;
  reg [31:0] _T_1696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3002;
  reg [31:0] _T_1696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3003;
  reg [31:0] _T_1697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3004;
  reg [31:0] _T_1697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3005;
  reg [31:0] _T_1698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3006;
  reg [31:0] _T_1698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3007;
  reg [31:0] _T_1699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3008;
  reg [31:0] _T_1699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3009;
  reg [31:0] _T_1702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3010;
  reg [31:0] _T_1702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3011;
  reg [31:0] _T_1703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3012;
  reg [31:0] _T_1703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3013;
  reg [31:0] _T_1704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3014;
  reg [31:0] _T_1704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3015;
  reg [31:0] _T_1705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3016;
  reg [31:0] _T_1705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3017;
  reg [31:0] _T_1706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3018;
  reg [31:0] _T_1706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3019;
  reg [31:0] _T_1707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3020;
  reg [31:0] _T_1707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3021;
  reg [31:0] _T_1708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3022;
  reg [31:0] _T_1708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3023;
  reg [31:0] _T_1709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3024;
  reg [31:0] _T_1709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3025;
  wire [31:0] _GEN_5042; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5043; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5044; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5045; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5046; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5047; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5050; // @[FFT.scala 35:12]
  wire [31:0] _GEN_5051; // @[FFT.scala 35:12]
  wire [31:0] _GEN_5052; // @[FFT.scala 35:12]
  wire [31:0] _GEN_5053; // @[FFT.scala 35:12]
  wire [31:0] _GEN_5054; // @[FFT.scala 35:12]
  wire [31:0] _GEN_5055; // @[FFT.scala 35:12]
  reg [31:0] _T_1715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3026;
  reg [31:0] _T_1715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3027;
  reg [31:0] _T_1716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3028;
  reg [31:0] _T_1716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3029;
  reg [31:0] _T_1717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3030;
  reg [31:0] _T_1717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3031;
  reg [31:0] _T_1718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3032;
  reg [31:0] _T_1718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3033;
  reg [31:0] _T_1719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3034;
  reg [31:0] _T_1719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3035;
  reg [31:0] _T_1720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3036;
  reg [31:0] _T_1720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3037;
  reg [31:0] _T_1721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3038;
  reg [31:0] _T_1721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3039;
  reg [31:0] _T_1722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3040;
  reg [31:0] _T_1722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3041;
  reg [31:0] _T_1725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3042;
  reg [31:0] _T_1725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3043;
  reg [31:0] _T_1726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3044;
  reg [31:0] _T_1726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3045;
  reg [31:0] _T_1727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3046;
  reg [31:0] _T_1727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3047;
  reg [31:0] _T_1728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3048;
  reg [31:0] _T_1728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3049;
  wire [31:0] _GEN_5082; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5083; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5086; // @[FFT.scala 35:12]
  wire [31:0] _GEN_5087; // @[FFT.scala 35:12]
  reg [31:0] _T_1734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3050;
  reg [31:0] _T_1734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3051;
  reg [31:0] _T_1735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3052;
  reg [31:0] _T_1735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3053;
  reg [31:0] _T_1736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3054;
  reg [31:0] _T_1736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3055;
  reg [31:0] _T_1737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3056;
  reg [31:0] _T_1737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3057;
  reg [31:0] _T_1740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3058;
  reg [31:0] _T_1740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3059;
  reg [31:0] _T_1741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3060;
  reg [31:0] _T_1741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3061;
  reg [31:0] _T_1747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3062;
  reg [31:0] _T_1747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3063;
  reg [31:0] _T_1748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3064;
  reg [31:0] _T_1748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3065;
  reg [31:0] _T_1751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3066;
  reg [31:0] _T_1751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3067;
  reg [31:0] out1D1_re; // @[FFT.scala 81:23]
  reg [31:0] _RAND_3068;
  reg [31:0] out1D1_im; // @[FFT.scala 81:23]
  reg [31:0] _RAND_3069;
  reg [31:0] _T_1752_re; // @[FFT.scala 85:22]
  reg [31:0] _RAND_3070;
  reg [31:0] _T_1752_im; // @[FFT.scala 85:22]
  reg [31:0] _RAND_3071;
  reg [31:0] _T_1753_re; // @[FFT.scala 86:22]
  reg [31:0] _RAND_3072;
  reg [31:0] _T_1753_im; // @[FFT.scala 86:22]
  reg [31:0] _RAND_3073;
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  Butterfly Butterfly_8 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_8_io_in1_re),
    .io_in1_im(Butterfly_8_io_in1_im),
    .io_in2_re(Butterfly_8_io_in2_re),
    .io_in2_im(Butterfly_8_io_in2_im),
    .io_wn_re(Butterfly_8_io_wn_re),
    .io_wn_im(Butterfly_8_io_wn_im),
    .io_out1_re(Butterfly_8_io_out1_re),
    .io_out1_im(Butterfly_8_io_out1_im),
    .io_out2_re(Butterfly_8_io_out2_re),
    .io_out2_im(Butterfly_8_io_out2_im)
  );
  Switch Switch_8 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_8_io_in1_re),
    .io_in1_im(Switch_8_io_in1_im),
    .io_in2_re(Switch_8_io_in2_re),
    .io_in2_im(Switch_8_io_in2_im),
    .io_sel(Switch_8_io_sel),
    .io_out1_re(Switch_8_io_out1_re),
    .io_out1_im(Switch_8_io_out1_im),
    .io_out2_re(Switch_8_io_out2_re),
    .io_out2_im(Switch_8_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign _T_1 = cnt + 10'h1; // @[FFT.scala 42:16]
  assign _GEN_2 = 9'h1 == cnt[8:0] ? $signed(32'shffff) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_3 = 9'h2 == cnt[8:0] ? $signed(32'shfffb) : $signed(_GEN_2); // @[FFT.scala 34:12]
  assign _GEN_4 = 9'h3 == cnt[8:0] ? $signed(32'shfff5) : $signed(_GEN_3); // @[FFT.scala 34:12]
  assign _GEN_5 = 9'h4 == cnt[8:0] ? $signed(32'shffec) : $signed(_GEN_4); // @[FFT.scala 34:12]
  assign _GEN_6 = 9'h5 == cnt[8:0] ? $signed(32'shffe1) : $signed(_GEN_5); // @[FFT.scala 34:12]
  assign _GEN_7 = 9'h6 == cnt[8:0] ? $signed(32'shffd4) : $signed(_GEN_6); // @[FFT.scala 34:12]
  assign _GEN_8 = 9'h7 == cnt[8:0] ? $signed(32'shffc4) : $signed(_GEN_7); // @[FFT.scala 34:12]
  assign _GEN_9 = 9'h8 == cnt[8:0] ? $signed(32'shffb1) : $signed(_GEN_8); // @[FFT.scala 34:12]
  assign _GEN_10 = 9'h9 == cnt[8:0] ? $signed(32'shff9c) : $signed(_GEN_9); // @[FFT.scala 34:12]
  assign _GEN_11 = 9'ha == cnt[8:0] ? $signed(32'shff85) : $signed(_GEN_10); // @[FFT.scala 34:12]
  assign _GEN_12 = 9'hb == cnt[8:0] ? $signed(32'shff6b) : $signed(_GEN_11); // @[FFT.scala 34:12]
  assign _GEN_13 = 9'hc == cnt[8:0] ? $signed(32'shff4e) : $signed(_GEN_12); // @[FFT.scala 34:12]
  assign _GEN_14 = 9'hd == cnt[8:0] ? $signed(32'shff30) : $signed(_GEN_13); // @[FFT.scala 34:12]
  assign _GEN_15 = 9'he == cnt[8:0] ? $signed(32'shff0e) : $signed(_GEN_14); // @[FFT.scala 34:12]
  assign _GEN_16 = 9'hf == cnt[8:0] ? $signed(32'shfeeb) : $signed(_GEN_15); // @[FFT.scala 34:12]
  assign _GEN_17 = 9'h10 == cnt[8:0] ? $signed(32'shfec4) : $signed(_GEN_16); // @[FFT.scala 34:12]
  assign _GEN_18 = 9'h11 == cnt[8:0] ? $signed(32'shfe9c) : $signed(_GEN_17); // @[FFT.scala 34:12]
  assign _GEN_19 = 9'h12 == cnt[8:0] ? $signed(32'shfe71) : $signed(_GEN_18); // @[FFT.scala 34:12]
  assign _GEN_20 = 9'h13 == cnt[8:0] ? $signed(32'shfe43) : $signed(_GEN_19); // @[FFT.scala 34:12]
  assign _GEN_21 = 9'h14 == cnt[8:0] ? $signed(32'shfe13) : $signed(_GEN_20); // @[FFT.scala 34:12]
  assign _GEN_22 = 9'h15 == cnt[8:0] ? $signed(32'shfde1) : $signed(_GEN_21); // @[FFT.scala 34:12]
  assign _GEN_23 = 9'h16 == cnt[8:0] ? $signed(32'shfdac) : $signed(_GEN_22); // @[FFT.scala 34:12]
  assign _GEN_24 = 9'h17 == cnt[8:0] ? $signed(32'shfd74) : $signed(_GEN_23); // @[FFT.scala 34:12]
  assign _GEN_25 = 9'h18 == cnt[8:0] ? $signed(32'shfd3b) : $signed(_GEN_24); // @[FFT.scala 34:12]
  assign _GEN_26 = 9'h19 == cnt[8:0] ? $signed(32'shfcfe) : $signed(_GEN_25); // @[FFT.scala 34:12]
  assign _GEN_27 = 9'h1a == cnt[8:0] ? $signed(32'shfcc0) : $signed(_GEN_26); // @[FFT.scala 34:12]
  assign _GEN_28 = 9'h1b == cnt[8:0] ? $signed(32'shfc7f) : $signed(_GEN_27); // @[FFT.scala 34:12]
  assign _GEN_29 = 9'h1c == cnt[8:0] ? $signed(32'shfc3b) : $signed(_GEN_28); // @[FFT.scala 34:12]
  assign _GEN_30 = 9'h1d == cnt[8:0] ? $signed(32'shfbf5) : $signed(_GEN_29); // @[FFT.scala 34:12]
  assign _GEN_31 = 9'h1e == cnt[8:0] ? $signed(32'shfbad) : $signed(_GEN_30); // @[FFT.scala 34:12]
  assign _GEN_32 = 9'h1f == cnt[8:0] ? $signed(32'shfb62) : $signed(_GEN_31); // @[FFT.scala 34:12]
  assign _GEN_33 = 9'h20 == cnt[8:0] ? $signed(32'shfb15) : $signed(_GEN_32); // @[FFT.scala 34:12]
  assign _GEN_34 = 9'h21 == cnt[8:0] ? $signed(32'shfac5) : $signed(_GEN_33); // @[FFT.scala 34:12]
  assign _GEN_35 = 9'h22 == cnt[8:0] ? $signed(32'shfa73) : $signed(_GEN_34); // @[FFT.scala 34:12]
  assign _GEN_36 = 9'h23 == cnt[8:0] ? $signed(32'shfa1f) : $signed(_GEN_35); // @[FFT.scala 34:12]
  assign _GEN_37 = 9'h24 == cnt[8:0] ? $signed(32'shf9c8) : $signed(_GEN_36); // @[FFT.scala 34:12]
  assign _GEN_38 = 9'h25 == cnt[8:0] ? $signed(32'shf96e) : $signed(_GEN_37); // @[FFT.scala 34:12]
  assign _GEN_39 = 9'h26 == cnt[8:0] ? $signed(32'shf913) : $signed(_GEN_38); // @[FFT.scala 34:12]
  assign _GEN_40 = 9'h27 == cnt[8:0] ? $signed(32'shf8b4) : $signed(_GEN_39); // @[FFT.scala 34:12]
  assign _GEN_41 = 9'h28 == cnt[8:0] ? $signed(32'shf854) : $signed(_GEN_40); // @[FFT.scala 34:12]
  assign _GEN_42 = 9'h29 == cnt[8:0] ? $signed(32'shf7f1) : $signed(_GEN_41); // @[FFT.scala 34:12]
  assign _GEN_43 = 9'h2a == cnt[8:0] ? $signed(32'shf78c) : $signed(_GEN_42); // @[FFT.scala 34:12]
  assign _GEN_44 = 9'h2b == cnt[8:0] ? $signed(32'shf724) : $signed(_GEN_43); // @[FFT.scala 34:12]
  assign _GEN_45 = 9'h2c == cnt[8:0] ? $signed(32'shf6ba) : $signed(_GEN_44); // @[FFT.scala 34:12]
  assign _GEN_46 = 9'h2d == cnt[8:0] ? $signed(32'shf64e) : $signed(_GEN_45); // @[FFT.scala 34:12]
  assign _GEN_47 = 9'h2e == cnt[8:0] ? $signed(32'shf5df) : $signed(_GEN_46); // @[FFT.scala 34:12]
  assign _GEN_48 = 9'h2f == cnt[8:0] ? $signed(32'shf56e) : $signed(_GEN_47); // @[FFT.scala 34:12]
  assign _GEN_49 = 9'h30 == cnt[8:0] ? $signed(32'shf4fa) : $signed(_GEN_48); // @[FFT.scala 34:12]
  assign _GEN_50 = 9'h31 == cnt[8:0] ? $signed(32'shf484) : $signed(_GEN_49); // @[FFT.scala 34:12]
  assign _GEN_51 = 9'h32 == cnt[8:0] ? $signed(32'shf40c) : $signed(_GEN_50); // @[FFT.scala 34:12]
  assign _GEN_52 = 9'h33 == cnt[8:0] ? $signed(32'shf391) : $signed(_GEN_51); // @[FFT.scala 34:12]
  assign _GEN_53 = 9'h34 == cnt[8:0] ? $signed(32'shf314) : $signed(_GEN_52); // @[FFT.scala 34:12]
  assign _GEN_54 = 9'h35 == cnt[8:0] ? $signed(32'shf295) : $signed(_GEN_53); // @[FFT.scala 34:12]
  assign _GEN_55 = 9'h36 == cnt[8:0] ? $signed(32'shf213) : $signed(_GEN_54); // @[FFT.scala 34:12]
  assign _GEN_56 = 9'h37 == cnt[8:0] ? $signed(32'shf18f) : $signed(_GEN_55); // @[FFT.scala 34:12]
  assign _GEN_57 = 9'h38 == cnt[8:0] ? $signed(32'shf109) : $signed(_GEN_56); // @[FFT.scala 34:12]
  assign _GEN_58 = 9'h39 == cnt[8:0] ? $signed(32'shf080) : $signed(_GEN_57); // @[FFT.scala 34:12]
  assign _GEN_59 = 9'h3a == cnt[8:0] ? $signed(32'sheff5) : $signed(_GEN_58); // @[FFT.scala 34:12]
  assign _GEN_60 = 9'h3b == cnt[8:0] ? $signed(32'shef68) : $signed(_GEN_59); // @[FFT.scala 34:12]
  assign _GEN_61 = 9'h3c == cnt[8:0] ? $signed(32'sheed9) : $signed(_GEN_60); // @[FFT.scala 34:12]
  assign _GEN_62 = 9'h3d == cnt[8:0] ? $signed(32'shee47) : $signed(_GEN_61); // @[FFT.scala 34:12]
  assign _GEN_63 = 9'h3e == cnt[8:0] ? $signed(32'shedb3) : $signed(_GEN_62); // @[FFT.scala 34:12]
  assign _GEN_64 = 9'h3f == cnt[8:0] ? $signed(32'shed1c) : $signed(_GEN_63); // @[FFT.scala 34:12]
  assign _GEN_65 = 9'h40 == cnt[8:0] ? $signed(32'shec83) : $signed(_GEN_64); // @[FFT.scala 34:12]
  assign _GEN_66 = 9'h41 == cnt[8:0] ? $signed(32'shebe8) : $signed(_GEN_65); // @[FFT.scala 34:12]
  assign _GEN_67 = 9'h42 == cnt[8:0] ? $signed(32'sheb4b) : $signed(_GEN_66); // @[FFT.scala 34:12]
  assign _GEN_68 = 9'h43 == cnt[8:0] ? $signed(32'sheaab) : $signed(_GEN_67); // @[FFT.scala 34:12]
  assign _GEN_69 = 9'h44 == cnt[8:0] ? $signed(32'shea0a) : $signed(_GEN_68); // @[FFT.scala 34:12]
  assign _GEN_70 = 9'h45 == cnt[8:0] ? $signed(32'she966) : $signed(_GEN_69); // @[FFT.scala 34:12]
  assign _GEN_71 = 9'h46 == cnt[8:0] ? $signed(32'she8bf) : $signed(_GEN_70); // @[FFT.scala 34:12]
  assign _GEN_72 = 9'h47 == cnt[8:0] ? $signed(32'she817) : $signed(_GEN_71); // @[FFT.scala 34:12]
  assign _GEN_73 = 9'h48 == cnt[8:0] ? $signed(32'she76c) : $signed(_GEN_72); // @[FFT.scala 34:12]
  assign _GEN_74 = 9'h49 == cnt[8:0] ? $signed(32'she6bf) : $signed(_GEN_73); // @[FFT.scala 34:12]
  assign _GEN_75 = 9'h4a == cnt[8:0] ? $signed(32'she610) : $signed(_GEN_74); // @[FFT.scala 34:12]
  assign _GEN_76 = 9'h4b == cnt[8:0] ? $signed(32'she55e) : $signed(_GEN_75); // @[FFT.scala 34:12]
  assign _GEN_77 = 9'h4c == cnt[8:0] ? $signed(32'she4aa) : $signed(_GEN_76); // @[FFT.scala 34:12]
  assign _GEN_78 = 9'h4d == cnt[8:0] ? $signed(32'she3f4) : $signed(_GEN_77); // @[FFT.scala 34:12]
  assign _GEN_79 = 9'h4e == cnt[8:0] ? $signed(32'she33c) : $signed(_GEN_78); // @[FFT.scala 34:12]
  assign _GEN_80 = 9'h4f == cnt[8:0] ? $signed(32'she282) : $signed(_GEN_79); // @[FFT.scala 34:12]
  assign _GEN_81 = 9'h50 == cnt[8:0] ? $signed(32'she1c6) : $signed(_GEN_80); // @[FFT.scala 34:12]
  assign _GEN_82 = 9'h51 == cnt[8:0] ? $signed(32'she107) : $signed(_GEN_81); // @[FFT.scala 34:12]
  assign _GEN_83 = 9'h52 == cnt[8:0] ? $signed(32'she046) : $signed(_GEN_82); // @[FFT.scala 34:12]
  assign _GEN_84 = 9'h53 == cnt[8:0] ? $signed(32'shdf83) : $signed(_GEN_83); // @[FFT.scala 34:12]
  assign _GEN_85 = 9'h54 == cnt[8:0] ? $signed(32'shdebe) : $signed(_GEN_84); // @[FFT.scala 34:12]
  assign _GEN_86 = 9'h55 == cnt[8:0] ? $signed(32'shddf7) : $signed(_GEN_85); // @[FFT.scala 34:12]
  assign _GEN_87 = 9'h56 == cnt[8:0] ? $signed(32'shdd2d) : $signed(_GEN_86); // @[FFT.scala 34:12]
  assign _GEN_88 = 9'h57 == cnt[8:0] ? $signed(32'shdc62) : $signed(_GEN_87); // @[FFT.scala 34:12]
  assign _GEN_89 = 9'h58 == cnt[8:0] ? $signed(32'shdb94) : $signed(_GEN_88); // @[FFT.scala 34:12]
  assign _GEN_90 = 9'h59 == cnt[8:0] ? $signed(32'shdac4) : $signed(_GEN_89); // @[FFT.scala 34:12]
  assign _GEN_91 = 9'h5a == cnt[8:0] ? $signed(32'shd9f2) : $signed(_GEN_90); // @[FFT.scala 34:12]
  assign _GEN_92 = 9'h5b == cnt[8:0] ? $signed(32'shd91e) : $signed(_GEN_91); // @[FFT.scala 34:12]
  assign _GEN_93 = 9'h5c == cnt[8:0] ? $signed(32'shd848) : $signed(_GEN_92); // @[FFT.scala 34:12]
  assign _GEN_94 = 9'h5d == cnt[8:0] ? $signed(32'shd770) : $signed(_GEN_93); // @[FFT.scala 34:12]
  assign _GEN_95 = 9'h5e == cnt[8:0] ? $signed(32'shd696) : $signed(_GEN_94); // @[FFT.scala 34:12]
  assign _GEN_96 = 9'h5f == cnt[8:0] ? $signed(32'shd5ba) : $signed(_GEN_95); // @[FFT.scala 34:12]
  assign _GEN_97 = 9'h60 == cnt[8:0] ? $signed(32'shd4db) : $signed(_GEN_96); // @[FFT.scala 34:12]
  assign _GEN_98 = 9'h61 == cnt[8:0] ? $signed(32'shd3fb) : $signed(_GEN_97); // @[FFT.scala 34:12]
  assign _GEN_99 = 9'h62 == cnt[8:0] ? $signed(32'shd318) : $signed(_GEN_98); // @[FFT.scala 34:12]
  assign _GEN_100 = 9'h63 == cnt[8:0] ? $signed(32'shd234) : $signed(_GEN_99); // @[FFT.scala 34:12]
  assign _GEN_101 = 9'h64 == cnt[8:0] ? $signed(32'shd14d) : $signed(_GEN_100); // @[FFT.scala 34:12]
  assign _GEN_102 = 9'h65 == cnt[8:0] ? $signed(32'shd065) : $signed(_GEN_101); // @[FFT.scala 34:12]
  assign _GEN_103 = 9'h66 == cnt[8:0] ? $signed(32'shcf7a) : $signed(_GEN_102); // @[FFT.scala 34:12]
  assign _GEN_104 = 9'h67 == cnt[8:0] ? $signed(32'shce8e) : $signed(_GEN_103); // @[FFT.scala 34:12]
  assign _GEN_105 = 9'h68 == cnt[8:0] ? $signed(32'shcd9f) : $signed(_GEN_104); // @[FFT.scala 34:12]
  assign _GEN_106 = 9'h69 == cnt[8:0] ? $signed(32'shccae) : $signed(_GEN_105); // @[FFT.scala 34:12]
  assign _GEN_107 = 9'h6a == cnt[8:0] ? $signed(32'shcbbc) : $signed(_GEN_106); // @[FFT.scala 34:12]
  assign _GEN_108 = 9'h6b == cnt[8:0] ? $signed(32'shcac7) : $signed(_GEN_107); // @[FFT.scala 34:12]
  assign _GEN_109 = 9'h6c == cnt[8:0] ? $signed(32'shc9d1) : $signed(_GEN_108); // @[FFT.scala 34:12]
  assign _GEN_110 = 9'h6d == cnt[8:0] ? $signed(32'shc8d9) : $signed(_GEN_109); // @[FFT.scala 34:12]
  assign _GEN_111 = 9'h6e == cnt[8:0] ? $signed(32'shc7de) : $signed(_GEN_110); // @[FFT.scala 34:12]
  assign _GEN_112 = 9'h6f == cnt[8:0] ? $signed(32'shc6e2) : $signed(_GEN_111); // @[FFT.scala 34:12]
  assign _GEN_113 = 9'h70 == cnt[8:0] ? $signed(32'shc5e4) : $signed(_GEN_112); // @[FFT.scala 34:12]
  assign _GEN_114 = 9'h71 == cnt[8:0] ? $signed(32'shc4e4) : $signed(_GEN_113); // @[FFT.scala 34:12]
  assign _GEN_115 = 9'h72 == cnt[8:0] ? $signed(32'shc3e2) : $signed(_GEN_114); // @[FFT.scala 34:12]
  assign _GEN_116 = 9'h73 == cnt[8:0] ? $signed(32'shc2de) : $signed(_GEN_115); // @[FFT.scala 34:12]
  assign _GEN_117 = 9'h74 == cnt[8:0] ? $signed(32'shc1d8) : $signed(_GEN_116); // @[FFT.scala 34:12]
  assign _GEN_118 = 9'h75 == cnt[8:0] ? $signed(32'shc0d1) : $signed(_GEN_117); // @[FFT.scala 34:12]
  assign _GEN_119 = 9'h76 == cnt[8:0] ? $signed(32'shbfc7) : $signed(_GEN_118); // @[FFT.scala 34:12]
  assign _GEN_120 = 9'h77 == cnt[8:0] ? $signed(32'shbebc) : $signed(_GEN_119); // @[FFT.scala 34:12]
  assign _GEN_121 = 9'h78 == cnt[8:0] ? $signed(32'shbdaf) : $signed(_GEN_120); // @[FFT.scala 34:12]
  assign _GEN_122 = 9'h79 == cnt[8:0] ? $signed(32'shbca0) : $signed(_GEN_121); // @[FFT.scala 34:12]
  assign _GEN_123 = 9'h7a == cnt[8:0] ? $signed(32'shbb8f) : $signed(_GEN_122); // @[FFT.scala 34:12]
  assign _GEN_124 = 9'h7b == cnt[8:0] ? $signed(32'shba7d) : $signed(_GEN_123); // @[FFT.scala 34:12]
  assign _GEN_125 = 9'h7c == cnt[8:0] ? $signed(32'shb968) : $signed(_GEN_124); // @[FFT.scala 34:12]
  assign _GEN_126 = 9'h7d == cnt[8:0] ? $signed(32'shb852) : $signed(_GEN_125); // @[FFT.scala 34:12]
  assign _GEN_127 = 9'h7e == cnt[8:0] ? $signed(32'shb73a) : $signed(_GEN_126); // @[FFT.scala 34:12]
  assign _GEN_128 = 9'h7f == cnt[8:0] ? $signed(32'shb620) : $signed(_GEN_127); // @[FFT.scala 34:12]
  assign _GEN_129 = 9'h80 == cnt[8:0] ? $signed(32'shb505) : $signed(_GEN_128); // @[FFT.scala 34:12]
  assign _GEN_130 = 9'h81 == cnt[8:0] ? $signed(32'shb3e8) : $signed(_GEN_129); // @[FFT.scala 34:12]
  assign _GEN_131 = 9'h82 == cnt[8:0] ? $signed(32'shb2c9) : $signed(_GEN_130); // @[FFT.scala 34:12]
  assign _GEN_132 = 9'h83 == cnt[8:0] ? $signed(32'shb1a8) : $signed(_GEN_131); // @[FFT.scala 34:12]
  assign _GEN_133 = 9'h84 == cnt[8:0] ? $signed(32'shb086) : $signed(_GEN_132); // @[FFT.scala 34:12]
  assign _GEN_134 = 9'h85 == cnt[8:0] ? $signed(32'shaf62) : $signed(_GEN_133); // @[FFT.scala 34:12]
  assign _GEN_135 = 9'h86 == cnt[8:0] ? $signed(32'shae3c) : $signed(_GEN_134); // @[FFT.scala 34:12]
  assign _GEN_136 = 9'h87 == cnt[8:0] ? $signed(32'shad14) : $signed(_GEN_135); // @[FFT.scala 34:12]
  assign _GEN_137 = 9'h88 == cnt[8:0] ? $signed(32'shabeb) : $signed(_GEN_136); // @[FFT.scala 34:12]
  assign _GEN_138 = 9'h89 == cnt[8:0] ? $signed(32'shaac1) : $signed(_GEN_137); // @[FFT.scala 34:12]
  assign _GEN_139 = 9'h8a == cnt[8:0] ? $signed(32'sha994) : $signed(_GEN_138); // @[FFT.scala 34:12]
  assign _GEN_140 = 9'h8b == cnt[8:0] ? $signed(32'sha866) : $signed(_GEN_139); // @[FFT.scala 34:12]
  assign _GEN_141 = 9'h8c == cnt[8:0] ? $signed(32'sha736) : $signed(_GEN_140); // @[FFT.scala 34:12]
  assign _GEN_142 = 9'h8d == cnt[8:0] ? $signed(32'sha605) : $signed(_GEN_141); // @[FFT.scala 34:12]
  assign _GEN_143 = 9'h8e == cnt[8:0] ? $signed(32'sha4d2) : $signed(_GEN_142); // @[FFT.scala 34:12]
  assign _GEN_144 = 9'h8f == cnt[8:0] ? $signed(32'sha39e) : $signed(_GEN_143); // @[FFT.scala 34:12]
  assign _GEN_145 = 9'h90 == cnt[8:0] ? $signed(32'sha268) : $signed(_GEN_144); // @[FFT.scala 34:12]
  assign _GEN_146 = 9'h91 == cnt[8:0] ? $signed(32'sha130) : $signed(_GEN_145); // @[FFT.scala 34:12]
  assign _GEN_147 = 9'h92 == cnt[8:0] ? $signed(32'sh9ff7) : $signed(_GEN_146); // @[FFT.scala 34:12]
  assign _GEN_148 = 9'h93 == cnt[8:0] ? $signed(32'sh9ebc) : $signed(_GEN_147); // @[FFT.scala 34:12]
  assign _GEN_149 = 9'h94 == cnt[8:0] ? $signed(32'sh9d80) : $signed(_GEN_148); // @[FFT.scala 34:12]
  assign _GEN_150 = 9'h95 == cnt[8:0] ? $signed(32'sh9c42) : $signed(_GEN_149); // @[FFT.scala 34:12]
  assign _GEN_151 = 9'h96 == cnt[8:0] ? $signed(32'sh9b03) : $signed(_GEN_150); // @[FFT.scala 34:12]
  assign _GEN_152 = 9'h97 == cnt[8:0] ? $signed(32'sh99c2) : $signed(_GEN_151); // @[FFT.scala 34:12]
  assign _GEN_153 = 9'h98 == cnt[8:0] ? $signed(32'sh9880) : $signed(_GEN_152); // @[FFT.scala 34:12]
  assign _GEN_154 = 9'h99 == cnt[8:0] ? $signed(32'sh973c) : $signed(_GEN_153); // @[FFT.scala 34:12]
  assign _GEN_155 = 9'h9a == cnt[8:0] ? $signed(32'sh95f7) : $signed(_GEN_154); // @[FFT.scala 34:12]
  assign _GEN_156 = 9'h9b == cnt[8:0] ? $signed(32'sh94b0) : $signed(_GEN_155); // @[FFT.scala 34:12]
  assign _GEN_157 = 9'h9c == cnt[8:0] ? $signed(32'sh9368) : $signed(_GEN_156); // @[FFT.scala 34:12]
  assign _GEN_158 = 9'h9d == cnt[8:0] ? $signed(32'sh921f) : $signed(_GEN_157); // @[FFT.scala 34:12]
  assign _GEN_159 = 9'h9e == cnt[8:0] ? $signed(32'sh90d4) : $signed(_GEN_158); // @[FFT.scala 34:12]
  assign _GEN_160 = 9'h9f == cnt[8:0] ? $signed(32'sh8f88) : $signed(_GEN_159); // @[FFT.scala 34:12]
  assign _GEN_161 = 9'ha0 == cnt[8:0] ? $signed(32'sh8e3a) : $signed(_GEN_160); // @[FFT.scala 34:12]
  assign _GEN_162 = 9'ha1 == cnt[8:0] ? $signed(32'sh8ceb) : $signed(_GEN_161); // @[FFT.scala 34:12]
  assign _GEN_163 = 9'ha2 == cnt[8:0] ? $signed(32'sh8b9a) : $signed(_GEN_162); // @[FFT.scala 34:12]
  assign _GEN_164 = 9'ha3 == cnt[8:0] ? $signed(32'sh8a49) : $signed(_GEN_163); // @[FFT.scala 34:12]
  assign _GEN_165 = 9'ha4 == cnt[8:0] ? $signed(32'sh88f6) : $signed(_GEN_164); // @[FFT.scala 34:12]
  assign _GEN_166 = 9'ha5 == cnt[8:0] ? $signed(32'sh87a1) : $signed(_GEN_165); // @[FFT.scala 34:12]
  assign _GEN_167 = 9'ha6 == cnt[8:0] ? $signed(32'sh864c) : $signed(_GEN_166); // @[FFT.scala 34:12]
  assign _GEN_168 = 9'ha7 == cnt[8:0] ? $signed(32'sh84f5) : $signed(_GEN_167); // @[FFT.scala 34:12]
  assign _GEN_169 = 9'ha8 == cnt[8:0] ? $signed(32'sh839c) : $signed(_GEN_168); // @[FFT.scala 34:12]
  assign _GEN_170 = 9'ha9 == cnt[8:0] ? $signed(32'sh8243) : $signed(_GEN_169); // @[FFT.scala 34:12]
  assign _GEN_171 = 9'haa == cnt[8:0] ? $signed(32'sh80e8) : $signed(_GEN_170); // @[FFT.scala 34:12]
  assign _GEN_172 = 9'hab == cnt[8:0] ? $signed(32'sh7f8c) : $signed(_GEN_171); // @[FFT.scala 34:12]
  assign _GEN_173 = 9'hac == cnt[8:0] ? $signed(32'sh7e2f) : $signed(_GEN_172); // @[FFT.scala 34:12]
  assign _GEN_174 = 9'had == cnt[8:0] ? $signed(32'sh7cd0) : $signed(_GEN_173); // @[FFT.scala 34:12]
  assign _GEN_175 = 9'hae == cnt[8:0] ? $signed(32'sh7b70) : $signed(_GEN_174); // @[FFT.scala 34:12]
  assign _GEN_176 = 9'haf == cnt[8:0] ? $signed(32'sh7a10) : $signed(_GEN_175); // @[FFT.scala 34:12]
  assign _GEN_177 = 9'hb0 == cnt[8:0] ? $signed(32'sh78ad) : $signed(_GEN_176); // @[FFT.scala 34:12]
  assign _GEN_178 = 9'hb1 == cnt[8:0] ? $signed(32'sh774a) : $signed(_GEN_177); // @[FFT.scala 34:12]
  assign _GEN_179 = 9'hb2 == cnt[8:0] ? $signed(32'sh75e6) : $signed(_GEN_178); // @[FFT.scala 34:12]
  assign _GEN_180 = 9'hb3 == cnt[8:0] ? $signed(32'sh7480) : $signed(_GEN_179); // @[FFT.scala 34:12]
  assign _GEN_181 = 9'hb4 == cnt[8:0] ? $signed(32'sh731a) : $signed(_GEN_180); // @[FFT.scala 34:12]
  assign _GEN_182 = 9'hb5 == cnt[8:0] ? $signed(32'sh71b2) : $signed(_GEN_181); // @[FFT.scala 34:12]
  assign _GEN_183 = 9'hb6 == cnt[8:0] ? $signed(32'sh7049) : $signed(_GEN_182); // @[FFT.scala 34:12]
  assign _GEN_184 = 9'hb7 == cnt[8:0] ? $signed(32'sh6edf) : $signed(_GEN_183); // @[FFT.scala 34:12]
  assign _GEN_185 = 9'hb8 == cnt[8:0] ? $signed(32'sh6d74) : $signed(_GEN_184); // @[FFT.scala 34:12]
  assign _GEN_186 = 9'hb9 == cnt[8:0] ? $signed(32'sh6c08) : $signed(_GEN_185); // @[FFT.scala 34:12]
  assign _GEN_187 = 9'hba == cnt[8:0] ? $signed(32'sh6a9b) : $signed(_GEN_186); // @[FFT.scala 34:12]
  assign _GEN_188 = 9'hbb == cnt[8:0] ? $signed(32'sh692d) : $signed(_GEN_187); // @[FFT.scala 34:12]
  assign _GEN_189 = 9'hbc == cnt[8:0] ? $signed(32'sh67be) : $signed(_GEN_188); // @[FFT.scala 34:12]
  assign _GEN_190 = 9'hbd == cnt[8:0] ? $signed(32'sh664e) : $signed(_GEN_189); // @[FFT.scala 34:12]
  assign _GEN_191 = 9'hbe == cnt[8:0] ? $signed(32'sh64dd) : $signed(_GEN_190); // @[FFT.scala 34:12]
  assign _GEN_192 = 9'hbf == cnt[8:0] ? $signed(32'sh636b) : $signed(_GEN_191); // @[FFT.scala 34:12]
  assign _GEN_193 = 9'hc0 == cnt[8:0] ? $signed(32'sh61f8) : $signed(_GEN_192); // @[FFT.scala 34:12]
  assign _GEN_194 = 9'hc1 == cnt[8:0] ? $signed(32'sh6084) : $signed(_GEN_193); // @[FFT.scala 34:12]
  assign _GEN_195 = 9'hc2 == cnt[8:0] ? $signed(32'sh5f0f) : $signed(_GEN_194); // @[FFT.scala 34:12]
  assign _GEN_196 = 9'hc3 == cnt[8:0] ? $signed(32'sh5d99) : $signed(_GEN_195); // @[FFT.scala 34:12]
  assign _GEN_197 = 9'hc4 == cnt[8:0] ? $signed(32'sh5c22) : $signed(_GEN_196); // @[FFT.scala 34:12]
  assign _GEN_198 = 9'hc5 == cnt[8:0] ? $signed(32'sh5aaa) : $signed(_GEN_197); // @[FFT.scala 34:12]
  assign _GEN_199 = 9'hc6 == cnt[8:0] ? $signed(32'sh5932) : $signed(_GEN_198); // @[FFT.scala 34:12]
  assign _GEN_200 = 9'hc7 == cnt[8:0] ? $signed(32'sh57b9) : $signed(_GEN_199); // @[FFT.scala 34:12]
  assign _GEN_201 = 9'hc8 == cnt[8:0] ? $signed(32'sh563e) : $signed(_GEN_200); // @[FFT.scala 34:12]
  assign _GEN_202 = 9'hc9 == cnt[8:0] ? $signed(32'sh54c3) : $signed(_GEN_201); // @[FFT.scala 34:12]
  assign _GEN_203 = 9'hca == cnt[8:0] ? $signed(32'sh5348) : $signed(_GEN_202); // @[FFT.scala 34:12]
  assign _GEN_204 = 9'hcb == cnt[8:0] ? $signed(32'sh51cb) : $signed(_GEN_203); // @[FFT.scala 34:12]
  assign _GEN_205 = 9'hcc == cnt[8:0] ? $signed(32'sh504d) : $signed(_GEN_204); // @[FFT.scala 34:12]
  assign _GEN_206 = 9'hcd == cnt[8:0] ? $signed(32'sh4ecf) : $signed(_GEN_205); // @[FFT.scala 34:12]
  assign _GEN_207 = 9'hce == cnt[8:0] ? $signed(32'sh4d50) : $signed(_GEN_206); // @[FFT.scala 34:12]
  assign _GEN_208 = 9'hcf == cnt[8:0] ? $signed(32'sh4bd1) : $signed(_GEN_207); // @[FFT.scala 34:12]
  assign _GEN_209 = 9'hd0 == cnt[8:0] ? $signed(32'sh4a50) : $signed(_GEN_208); // @[FFT.scala 34:12]
  assign _GEN_210 = 9'hd1 == cnt[8:0] ? $signed(32'sh48cf) : $signed(_GEN_209); // @[FFT.scala 34:12]
  assign _GEN_211 = 9'hd2 == cnt[8:0] ? $signed(32'sh474d) : $signed(_GEN_210); // @[FFT.scala 34:12]
  assign _GEN_212 = 9'hd3 == cnt[8:0] ? $signed(32'sh45cb) : $signed(_GEN_211); // @[FFT.scala 34:12]
  assign _GEN_213 = 9'hd4 == cnt[8:0] ? $signed(32'sh4447) : $signed(_GEN_212); // @[FFT.scala 34:12]
  assign _GEN_214 = 9'hd5 == cnt[8:0] ? $signed(32'sh42c3) : $signed(_GEN_213); // @[FFT.scala 34:12]
  assign _GEN_215 = 9'hd6 == cnt[8:0] ? $signed(32'sh413f) : $signed(_GEN_214); // @[FFT.scala 34:12]
  assign _GEN_216 = 9'hd7 == cnt[8:0] ? $signed(32'sh3fba) : $signed(_GEN_215); // @[FFT.scala 34:12]
  assign _GEN_217 = 9'hd8 == cnt[8:0] ? $signed(32'sh3e34) : $signed(_GEN_216); // @[FFT.scala 34:12]
  assign _GEN_218 = 9'hd9 == cnt[8:0] ? $signed(32'sh3cae) : $signed(_GEN_217); // @[FFT.scala 34:12]
  assign _GEN_219 = 9'hda == cnt[8:0] ? $signed(32'sh3b27) : $signed(_GEN_218); // @[FFT.scala 34:12]
  assign _GEN_220 = 9'hdb == cnt[8:0] ? $signed(32'sh399f) : $signed(_GEN_219); // @[FFT.scala 34:12]
  assign _GEN_221 = 9'hdc == cnt[8:0] ? $signed(32'sh3817) : $signed(_GEN_220); // @[FFT.scala 34:12]
  assign _GEN_222 = 9'hdd == cnt[8:0] ? $signed(32'sh368e) : $signed(_GEN_221); // @[FFT.scala 34:12]
  assign _GEN_223 = 9'hde == cnt[8:0] ? $signed(32'sh3505) : $signed(_GEN_222); // @[FFT.scala 34:12]
  assign _GEN_224 = 9'hdf == cnt[8:0] ? $signed(32'sh337c) : $signed(_GEN_223); // @[FFT.scala 34:12]
  assign _GEN_225 = 9'he0 == cnt[8:0] ? $signed(32'sh31f1) : $signed(_GEN_224); // @[FFT.scala 34:12]
  assign _GEN_226 = 9'he1 == cnt[8:0] ? $signed(32'sh3067) : $signed(_GEN_225); // @[FFT.scala 34:12]
  assign _GEN_227 = 9'he2 == cnt[8:0] ? $signed(32'sh2edc) : $signed(_GEN_226); // @[FFT.scala 34:12]
  assign _GEN_228 = 9'he3 == cnt[8:0] ? $signed(32'sh2d50) : $signed(_GEN_227); // @[FFT.scala 34:12]
  assign _GEN_229 = 9'he4 == cnt[8:0] ? $signed(32'sh2bc4) : $signed(_GEN_228); // @[FFT.scala 34:12]
  assign _GEN_230 = 9'he5 == cnt[8:0] ? $signed(32'sh2a38) : $signed(_GEN_229); // @[FFT.scala 34:12]
  assign _GEN_231 = 9'he6 == cnt[8:0] ? $signed(32'sh28ab) : $signed(_GEN_230); // @[FFT.scala 34:12]
  assign _GEN_232 = 9'he7 == cnt[8:0] ? $signed(32'sh271e) : $signed(_GEN_231); // @[FFT.scala 34:12]
  assign _GEN_233 = 9'he8 == cnt[8:0] ? $signed(32'sh2590) : $signed(_GEN_232); // @[FFT.scala 34:12]
  assign _GEN_234 = 9'he9 == cnt[8:0] ? $signed(32'sh2402) : $signed(_GEN_233); // @[FFT.scala 34:12]
  assign _GEN_235 = 9'hea == cnt[8:0] ? $signed(32'sh2274) : $signed(_GEN_234); // @[FFT.scala 34:12]
  assign _GEN_236 = 9'heb == cnt[8:0] ? $signed(32'sh20e5) : $signed(_GEN_235); // @[FFT.scala 34:12]
  assign _GEN_237 = 9'hec == cnt[8:0] ? $signed(32'sh1f56) : $signed(_GEN_236); // @[FFT.scala 34:12]
  assign _GEN_238 = 9'hed == cnt[8:0] ? $signed(32'sh1dc7) : $signed(_GEN_237); // @[FFT.scala 34:12]
  assign _GEN_239 = 9'hee == cnt[8:0] ? $signed(32'sh1c38) : $signed(_GEN_238); // @[FFT.scala 34:12]
  assign _GEN_240 = 9'hef == cnt[8:0] ? $signed(32'sh1aa8) : $signed(_GEN_239); // @[FFT.scala 34:12]
  assign _GEN_241 = 9'hf0 == cnt[8:0] ? $signed(32'sh1918) : $signed(_GEN_240); // @[FFT.scala 34:12]
  assign _GEN_242 = 9'hf1 == cnt[8:0] ? $signed(32'sh1787) : $signed(_GEN_241); // @[FFT.scala 34:12]
  assign _GEN_243 = 9'hf2 == cnt[8:0] ? $signed(32'sh15f7) : $signed(_GEN_242); // @[FFT.scala 34:12]
  assign _GEN_244 = 9'hf3 == cnt[8:0] ? $signed(32'sh1466) : $signed(_GEN_243); // @[FFT.scala 34:12]
  assign _GEN_245 = 9'hf4 == cnt[8:0] ? $signed(32'sh12d5) : $signed(_GEN_244); // @[FFT.scala 34:12]
  assign _GEN_246 = 9'hf5 == cnt[8:0] ? $signed(32'sh1144) : $signed(_GEN_245); // @[FFT.scala 34:12]
  assign _GEN_247 = 9'hf6 == cnt[8:0] ? $signed(32'shfb3) : $signed(_GEN_246); // @[FFT.scala 34:12]
  assign _GEN_248 = 9'hf7 == cnt[8:0] ? $signed(32'she21) : $signed(_GEN_247); // @[FFT.scala 34:12]
  assign _GEN_249 = 9'hf8 == cnt[8:0] ? $signed(32'shc90) : $signed(_GEN_248); // @[FFT.scala 34:12]
  assign _GEN_250 = 9'hf9 == cnt[8:0] ? $signed(32'shafe) : $signed(_GEN_249); // @[FFT.scala 34:12]
  assign _GEN_251 = 9'hfa == cnt[8:0] ? $signed(32'sh96c) : $signed(_GEN_250); // @[FFT.scala 34:12]
  assign _GEN_252 = 9'hfb == cnt[8:0] ? $signed(32'sh7da) : $signed(_GEN_251); // @[FFT.scala 34:12]
  assign _GEN_253 = 9'hfc == cnt[8:0] ? $signed(32'sh648) : $signed(_GEN_252); // @[FFT.scala 34:12]
  assign _GEN_254 = 9'hfd == cnt[8:0] ? $signed(32'sh4b6) : $signed(_GEN_253); // @[FFT.scala 34:12]
  assign _GEN_255 = 9'hfe == cnt[8:0] ? $signed(32'sh324) : $signed(_GEN_254); // @[FFT.scala 34:12]
  assign _GEN_256 = 9'hff == cnt[8:0] ? $signed(32'sh192) : $signed(_GEN_255); // @[FFT.scala 34:12]
  assign _GEN_257 = 9'h100 == cnt[8:0] ? $signed(32'sh0) : $signed(_GEN_256); // @[FFT.scala 34:12]
  assign _GEN_258 = 9'h101 == cnt[8:0] ? $signed(-32'sh192) : $signed(_GEN_257); // @[FFT.scala 34:12]
  assign _GEN_259 = 9'h102 == cnt[8:0] ? $signed(-32'sh324) : $signed(_GEN_258); // @[FFT.scala 34:12]
  assign _GEN_260 = 9'h103 == cnt[8:0] ? $signed(-32'sh4b6) : $signed(_GEN_259); // @[FFT.scala 34:12]
  assign _GEN_261 = 9'h104 == cnt[8:0] ? $signed(-32'sh648) : $signed(_GEN_260); // @[FFT.scala 34:12]
  assign _GEN_262 = 9'h105 == cnt[8:0] ? $signed(-32'sh7da) : $signed(_GEN_261); // @[FFT.scala 34:12]
  assign _GEN_263 = 9'h106 == cnt[8:0] ? $signed(-32'sh96c) : $signed(_GEN_262); // @[FFT.scala 34:12]
  assign _GEN_264 = 9'h107 == cnt[8:0] ? $signed(-32'shafe) : $signed(_GEN_263); // @[FFT.scala 34:12]
  assign _GEN_265 = 9'h108 == cnt[8:0] ? $signed(-32'shc90) : $signed(_GEN_264); // @[FFT.scala 34:12]
  assign _GEN_266 = 9'h109 == cnt[8:0] ? $signed(-32'she21) : $signed(_GEN_265); // @[FFT.scala 34:12]
  assign _GEN_267 = 9'h10a == cnt[8:0] ? $signed(-32'shfb3) : $signed(_GEN_266); // @[FFT.scala 34:12]
  assign _GEN_268 = 9'h10b == cnt[8:0] ? $signed(-32'sh1144) : $signed(_GEN_267); // @[FFT.scala 34:12]
  assign _GEN_269 = 9'h10c == cnt[8:0] ? $signed(-32'sh12d5) : $signed(_GEN_268); // @[FFT.scala 34:12]
  assign _GEN_270 = 9'h10d == cnt[8:0] ? $signed(-32'sh1466) : $signed(_GEN_269); // @[FFT.scala 34:12]
  assign _GEN_271 = 9'h10e == cnt[8:0] ? $signed(-32'sh15f7) : $signed(_GEN_270); // @[FFT.scala 34:12]
  assign _GEN_272 = 9'h10f == cnt[8:0] ? $signed(-32'sh1787) : $signed(_GEN_271); // @[FFT.scala 34:12]
  assign _GEN_273 = 9'h110 == cnt[8:0] ? $signed(-32'sh1918) : $signed(_GEN_272); // @[FFT.scala 34:12]
  assign _GEN_274 = 9'h111 == cnt[8:0] ? $signed(-32'sh1aa8) : $signed(_GEN_273); // @[FFT.scala 34:12]
  assign _GEN_275 = 9'h112 == cnt[8:0] ? $signed(-32'sh1c38) : $signed(_GEN_274); // @[FFT.scala 34:12]
  assign _GEN_276 = 9'h113 == cnt[8:0] ? $signed(-32'sh1dc7) : $signed(_GEN_275); // @[FFT.scala 34:12]
  assign _GEN_277 = 9'h114 == cnt[8:0] ? $signed(-32'sh1f56) : $signed(_GEN_276); // @[FFT.scala 34:12]
  assign _GEN_278 = 9'h115 == cnt[8:0] ? $signed(-32'sh20e5) : $signed(_GEN_277); // @[FFT.scala 34:12]
  assign _GEN_279 = 9'h116 == cnt[8:0] ? $signed(-32'sh2274) : $signed(_GEN_278); // @[FFT.scala 34:12]
  assign _GEN_280 = 9'h117 == cnt[8:0] ? $signed(-32'sh2402) : $signed(_GEN_279); // @[FFT.scala 34:12]
  assign _GEN_281 = 9'h118 == cnt[8:0] ? $signed(-32'sh2590) : $signed(_GEN_280); // @[FFT.scala 34:12]
  assign _GEN_282 = 9'h119 == cnt[8:0] ? $signed(-32'sh271e) : $signed(_GEN_281); // @[FFT.scala 34:12]
  assign _GEN_283 = 9'h11a == cnt[8:0] ? $signed(-32'sh28ab) : $signed(_GEN_282); // @[FFT.scala 34:12]
  assign _GEN_284 = 9'h11b == cnt[8:0] ? $signed(-32'sh2a38) : $signed(_GEN_283); // @[FFT.scala 34:12]
  assign _GEN_285 = 9'h11c == cnt[8:0] ? $signed(-32'sh2bc4) : $signed(_GEN_284); // @[FFT.scala 34:12]
  assign _GEN_286 = 9'h11d == cnt[8:0] ? $signed(-32'sh2d50) : $signed(_GEN_285); // @[FFT.scala 34:12]
  assign _GEN_287 = 9'h11e == cnt[8:0] ? $signed(-32'sh2edc) : $signed(_GEN_286); // @[FFT.scala 34:12]
  assign _GEN_288 = 9'h11f == cnt[8:0] ? $signed(-32'sh3067) : $signed(_GEN_287); // @[FFT.scala 34:12]
  assign _GEN_289 = 9'h120 == cnt[8:0] ? $signed(-32'sh31f1) : $signed(_GEN_288); // @[FFT.scala 34:12]
  assign _GEN_290 = 9'h121 == cnt[8:0] ? $signed(-32'sh337c) : $signed(_GEN_289); // @[FFT.scala 34:12]
  assign _GEN_291 = 9'h122 == cnt[8:0] ? $signed(-32'sh3505) : $signed(_GEN_290); // @[FFT.scala 34:12]
  assign _GEN_292 = 9'h123 == cnt[8:0] ? $signed(-32'sh368e) : $signed(_GEN_291); // @[FFT.scala 34:12]
  assign _GEN_293 = 9'h124 == cnt[8:0] ? $signed(-32'sh3817) : $signed(_GEN_292); // @[FFT.scala 34:12]
  assign _GEN_294 = 9'h125 == cnt[8:0] ? $signed(-32'sh399f) : $signed(_GEN_293); // @[FFT.scala 34:12]
  assign _GEN_295 = 9'h126 == cnt[8:0] ? $signed(-32'sh3b27) : $signed(_GEN_294); // @[FFT.scala 34:12]
  assign _GEN_296 = 9'h127 == cnt[8:0] ? $signed(-32'sh3cae) : $signed(_GEN_295); // @[FFT.scala 34:12]
  assign _GEN_297 = 9'h128 == cnt[8:0] ? $signed(-32'sh3e34) : $signed(_GEN_296); // @[FFT.scala 34:12]
  assign _GEN_298 = 9'h129 == cnt[8:0] ? $signed(-32'sh3fba) : $signed(_GEN_297); // @[FFT.scala 34:12]
  assign _GEN_299 = 9'h12a == cnt[8:0] ? $signed(-32'sh413f) : $signed(_GEN_298); // @[FFT.scala 34:12]
  assign _GEN_300 = 9'h12b == cnt[8:0] ? $signed(-32'sh42c3) : $signed(_GEN_299); // @[FFT.scala 34:12]
  assign _GEN_301 = 9'h12c == cnt[8:0] ? $signed(-32'sh4447) : $signed(_GEN_300); // @[FFT.scala 34:12]
  assign _GEN_302 = 9'h12d == cnt[8:0] ? $signed(-32'sh45cb) : $signed(_GEN_301); // @[FFT.scala 34:12]
  assign _GEN_303 = 9'h12e == cnt[8:0] ? $signed(-32'sh474d) : $signed(_GEN_302); // @[FFT.scala 34:12]
  assign _GEN_304 = 9'h12f == cnt[8:0] ? $signed(-32'sh48cf) : $signed(_GEN_303); // @[FFT.scala 34:12]
  assign _GEN_305 = 9'h130 == cnt[8:0] ? $signed(-32'sh4a50) : $signed(_GEN_304); // @[FFT.scala 34:12]
  assign _GEN_306 = 9'h131 == cnt[8:0] ? $signed(-32'sh4bd1) : $signed(_GEN_305); // @[FFT.scala 34:12]
  assign _GEN_307 = 9'h132 == cnt[8:0] ? $signed(-32'sh4d50) : $signed(_GEN_306); // @[FFT.scala 34:12]
  assign _GEN_308 = 9'h133 == cnt[8:0] ? $signed(-32'sh4ecf) : $signed(_GEN_307); // @[FFT.scala 34:12]
  assign _GEN_309 = 9'h134 == cnt[8:0] ? $signed(-32'sh504d) : $signed(_GEN_308); // @[FFT.scala 34:12]
  assign _GEN_310 = 9'h135 == cnt[8:0] ? $signed(-32'sh51cb) : $signed(_GEN_309); // @[FFT.scala 34:12]
  assign _GEN_311 = 9'h136 == cnt[8:0] ? $signed(-32'sh5348) : $signed(_GEN_310); // @[FFT.scala 34:12]
  assign _GEN_312 = 9'h137 == cnt[8:0] ? $signed(-32'sh54c3) : $signed(_GEN_311); // @[FFT.scala 34:12]
  assign _GEN_313 = 9'h138 == cnt[8:0] ? $signed(-32'sh563e) : $signed(_GEN_312); // @[FFT.scala 34:12]
  assign _GEN_314 = 9'h139 == cnt[8:0] ? $signed(-32'sh57b9) : $signed(_GEN_313); // @[FFT.scala 34:12]
  assign _GEN_315 = 9'h13a == cnt[8:0] ? $signed(-32'sh5932) : $signed(_GEN_314); // @[FFT.scala 34:12]
  assign _GEN_316 = 9'h13b == cnt[8:0] ? $signed(-32'sh5aaa) : $signed(_GEN_315); // @[FFT.scala 34:12]
  assign _GEN_317 = 9'h13c == cnt[8:0] ? $signed(-32'sh5c22) : $signed(_GEN_316); // @[FFT.scala 34:12]
  assign _GEN_318 = 9'h13d == cnt[8:0] ? $signed(-32'sh5d99) : $signed(_GEN_317); // @[FFT.scala 34:12]
  assign _GEN_319 = 9'h13e == cnt[8:0] ? $signed(-32'sh5f0f) : $signed(_GEN_318); // @[FFT.scala 34:12]
  assign _GEN_320 = 9'h13f == cnt[8:0] ? $signed(-32'sh6084) : $signed(_GEN_319); // @[FFT.scala 34:12]
  assign _GEN_321 = 9'h140 == cnt[8:0] ? $signed(-32'sh61f8) : $signed(_GEN_320); // @[FFT.scala 34:12]
  assign _GEN_322 = 9'h141 == cnt[8:0] ? $signed(-32'sh636b) : $signed(_GEN_321); // @[FFT.scala 34:12]
  assign _GEN_323 = 9'h142 == cnt[8:0] ? $signed(-32'sh64dd) : $signed(_GEN_322); // @[FFT.scala 34:12]
  assign _GEN_324 = 9'h143 == cnt[8:0] ? $signed(-32'sh664e) : $signed(_GEN_323); // @[FFT.scala 34:12]
  assign _GEN_325 = 9'h144 == cnt[8:0] ? $signed(-32'sh67be) : $signed(_GEN_324); // @[FFT.scala 34:12]
  assign _GEN_326 = 9'h145 == cnt[8:0] ? $signed(-32'sh692d) : $signed(_GEN_325); // @[FFT.scala 34:12]
  assign _GEN_327 = 9'h146 == cnt[8:0] ? $signed(-32'sh6a9b) : $signed(_GEN_326); // @[FFT.scala 34:12]
  assign _GEN_328 = 9'h147 == cnt[8:0] ? $signed(-32'sh6c08) : $signed(_GEN_327); // @[FFT.scala 34:12]
  assign _GEN_329 = 9'h148 == cnt[8:0] ? $signed(-32'sh6d74) : $signed(_GEN_328); // @[FFT.scala 34:12]
  assign _GEN_330 = 9'h149 == cnt[8:0] ? $signed(-32'sh6edf) : $signed(_GEN_329); // @[FFT.scala 34:12]
  assign _GEN_331 = 9'h14a == cnt[8:0] ? $signed(-32'sh7049) : $signed(_GEN_330); // @[FFT.scala 34:12]
  assign _GEN_332 = 9'h14b == cnt[8:0] ? $signed(-32'sh71b2) : $signed(_GEN_331); // @[FFT.scala 34:12]
  assign _GEN_333 = 9'h14c == cnt[8:0] ? $signed(-32'sh731a) : $signed(_GEN_332); // @[FFT.scala 34:12]
  assign _GEN_334 = 9'h14d == cnt[8:0] ? $signed(-32'sh7480) : $signed(_GEN_333); // @[FFT.scala 34:12]
  assign _GEN_335 = 9'h14e == cnt[8:0] ? $signed(-32'sh75e6) : $signed(_GEN_334); // @[FFT.scala 34:12]
  assign _GEN_336 = 9'h14f == cnt[8:0] ? $signed(-32'sh774a) : $signed(_GEN_335); // @[FFT.scala 34:12]
  assign _GEN_337 = 9'h150 == cnt[8:0] ? $signed(-32'sh78ad) : $signed(_GEN_336); // @[FFT.scala 34:12]
  assign _GEN_338 = 9'h151 == cnt[8:0] ? $signed(-32'sh7a10) : $signed(_GEN_337); // @[FFT.scala 34:12]
  assign _GEN_339 = 9'h152 == cnt[8:0] ? $signed(-32'sh7b70) : $signed(_GEN_338); // @[FFT.scala 34:12]
  assign _GEN_340 = 9'h153 == cnt[8:0] ? $signed(-32'sh7cd0) : $signed(_GEN_339); // @[FFT.scala 34:12]
  assign _GEN_341 = 9'h154 == cnt[8:0] ? $signed(-32'sh7e2f) : $signed(_GEN_340); // @[FFT.scala 34:12]
  assign _GEN_342 = 9'h155 == cnt[8:0] ? $signed(-32'sh7f8c) : $signed(_GEN_341); // @[FFT.scala 34:12]
  assign _GEN_343 = 9'h156 == cnt[8:0] ? $signed(-32'sh80e8) : $signed(_GEN_342); // @[FFT.scala 34:12]
  assign _GEN_344 = 9'h157 == cnt[8:0] ? $signed(-32'sh8243) : $signed(_GEN_343); // @[FFT.scala 34:12]
  assign _GEN_345 = 9'h158 == cnt[8:0] ? $signed(-32'sh839c) : $signed(_GEN_344); // @[FFT.scala 34:12]
  assign _GEN_346 = 9'h159 == cnt[8:0] ? $signed(-32'sh84f5) : $signed(_GEN_345); // @[FFT.scala 34:12]
  assign _GEN_347 = 9'h15a == cnt[8:0] ? $signed(-32'sh864c) : $signed(_GEN_346); // @[FFT.scala 34:12]
  assign _GEN_348 = 9'h15b == cnt[8:0] ? $signed(-32'sh87a1) : $signed(_GEN_347); // @[FFT.scala 34:12]
  assign _GEN_349 = 9'h15c == cnt[8:0] ? $signed(-32'sh88f6) : $signed(_GEN_348); // @[FFT.scala 34:12]
  assign _GEN_350 = 9'h15d == cnt[8:0] ? $signed(-32'sh8a49) : $signed(_GEN_349); // @[FFT.scala 34:12]
  assign _GEN_351 = 9'h15e == cnt[8:0] ? $signed(-32'sh8b9a) : $signed(_GEN_350); // @[FFT.scala 34:12]
  assign _GEN_352 = 9'h15f == cnt[8:0] ? $signed(-32'sh8ceb) : $signed(_GEN_351); // @[FFT.scala 34:12]
  assign _GEN_353 = 9'h160 == cnt[8:0] ? $signed(-32'sh8e3a) : $signed(_GEN_352); // @[FFT.scala 34:12]
  assign _GEN_354 = 9'h161 == cnt[8:0] ? $signed(-32'sh8f88) : $signed(_GEN_353); // @[FFT.scala 34:12]
  assign _GEN_355 = 9'h162 == cnt[8:0] ? $signed(-32'sh90d4) : $signed(_GEN_354); // @[FFT.scala 34:12]
  assign _GEN_356 = 9'h163 == cnt[8:0] ? $signed(-32'sh921f) : $signed(_GEN_355); // @[FFT.scala 34:12]
  assign _GEN_357 = 9'h164 == cnt[8:0] ? $signed(-32'sh9368) : $signed(_GEN_356); // @[FFT.scala 34:12]
  assign _GEN_358 = 9'h165 == cnt[8:0] ? $signed(-32'sh94b0) : $signed(_GEN_357); // @[FFT.scala 34:12]
  assign _GEN_359 = 9'h166 == cnt[8:0] ? $signed(-32'sh95f7) : $signed(_GEN_358); // @[FFT.scala 34:12]
  assign _GEN_360 = 9'h167 == cnt[8:0] ? $signed(-32'sh973c) : $signed(_GEN_359); // @[FFT.scala 34:12]
  assign _GEN_361 = 9'h168 == cnt[8:0] ? $signed(-32'sh9880) : $signed(_GEN_360); // @[FFT.scala 34:12]
  assign _GEN_362 = 9'h169 == cnt[8:0] ? $signed(-32'sh99c2) : $signed(_GEN_361); // @[FFT.scala 34:12]
  assign _GEN_363 = 9'h16a == cnt[8:0] ? $signed(-32'sh9b03) : $signed(_GEN_362); // @[FFT.scala 34:12]
  assign _GEN_364 = 9'h16b == cnt[8:0] ? $signed(-32'sh9c42) : $signed(_GEN_363); // @[FFT.scala 34:12]
  assign _GEN_365 = 9'h16c == cnt[8:0] ? $signed(-32'sh9d80) : $signed(_GEN_364); // @[FFT.scala 34:12]
  assign _GEN_366 = 9'h16d == cnt[8:0] ? $signed(-32'sh9ebc) : $signed(_GEN_365); // @[FFT.scala 34:12]
  assign _GEN_367 = 9'h16e == cnt[8:0] ? $signed(-32'sh9ff7) : $signed(_GEN_366); // @[FFT.scala 34:12]
  assign _GEN_368 = 9'h16f == cnt[8:0] ? $signed(-32'sha130) : $signed(_GEN_367); // @[FFT.scala 34:12]
  assign _GEN_369 = 9'h170 == cnt[8:0] ? $signed(-32'sha268) : $signed(_GEN_368); // @[FFT.scala 34:12]
  assign _GEN_370 = 9'h171 == cnt[8:0] ? $signed(-32'sha39e) : $signed(_GEN_369); // @[FFT.scala 34:12]
  assign _GEN_371 = 9'h172 == cnt[8:0] ? $signed(-32'sha4d2) : $signed(_GEN_370); // @[FFT.scala 34:12]
  assign _GEN_372 = 9'h173 == cnt[8:0] ? $signed(-32'sha605) : $signed(_GEN_371); // @[FFT.scala 34:12]
  assign _GEN_373 = 9'h174 == cnt[8:0] ? $signed(-32'sha736) : $signed(_GEN_372); // @[FFT.scala 34:12]
  assign _GEN_374 = 9'h175 == cnt[8:0] ? $signed(-32'sha866) : $signed(_GEN_373); // @[FFT.scala 34:12]
  assign _GEN_375 = 9'h176 == cnt[8:0] ? $signed(-32'sha994) : $signed(_GEN_374); // @[FFT.scala 34:12]
  assign _GEN_376 = 9'h177 == cnt[8:0] ? $signed(-32'shaac1) : $signed(_GEN_375); // @[FFT.scala 34:12]
  assign _GEN_377 = 9'h178 == cnt[8:0] ? $signed(-32'shabeb) : $signed(_GEN_376); // @[FFT.scala 34:12]
  assign _GEN_378 = 9'h179 == cnt[8:0] ? $signed(-32'shad14) : $signed(_GEN_377); // @[FFT.scala 34:12]
  assign _GEN_379 = 9'h17a == cnt[8:0] ? $signed(-32'shae3c) : $signed(_GEN_378); // @[FFT.scala 34:12]
  assign _GEN_380 = 9'h17b == cnt[8:0] ? $signed(-32'shaf62) : $signed(_GEN_379); // @[FFT.scala 34:12]
  assign _GEN_381 = 9'h17c == cnt[8:0] ? $signed(-32'shb086) : $signed(_GEN_380); // @[FFT.scala 34:12]
  assign _GEN_382 = 9'h17d == cnt[8:0] ? $signed(-32'shb1a8) : $signed(_GEN_381); // @[FFT.scala 34:12]
  assign _GEN_383 = 9'h17e == cnt[8:0] ? $signed(-32'shb2c9) : $signed(_GEN_382); // @[FFT.scala 34:12]
  assign _GEN_384 = 9'h17f == cnt[8:0] ? $signed(-32'shb3e8) : $signed(_GEN_383); // @[FFT.scala 34:12]
  assign _GEN_385 = 9'h180 == cnt[8:0] ? $signed(-32'shb505) : $signed(_GEN_384); // @[FFT.scala 34:12]
  assign _GEN_386 = 9'h181 == cnt[8:0] ? $signed(-32'shb620) : $signed(_GEN_385); // @[FFT.scala 34:12]
  assign _GEN_387 = 9'h182 == cnt[8:0] ? $signed(-32'shb73a) : $signed(_GEN_386); // @[FFT.scala 34:12]
  assign _GEN_388 = 9'h183 == cnt[8:0] ? $signed(-32'shb852) : $signed(_GEN_387); // @[FFT.scala 34:12]
  assign _GEN_389 = 9'h184 == cnt[8:0] ? $signed(-32'shb968) : $signed(_GEN_388); // @[FFT.scala 34:12]
  assign _GEN_390 = 9'h185 == cnt[8:0] ? $signed(-32'shba7d) : $signed(_GEN_389); // @[FFT.scala 34:12]
  assign _GEN_391 = 9'h186 == cnt[8:0] ? $signed(-32'shbb8f) : $signed(_GEN_390); // @[FFT.scala 34:12]
  assign _GEN_392 = 9'h187 == cnt[8:0] ? $signed(-32'shbca0) : $signed(_GEN_391); // @[FFT.scala 34:12]
  assign _GEN_393 = 9'h188 == cnt[8:0] ? $signed(-32'shbdaf) : $signed(_GEN_392); // @[FFT.scala 34:12]
  assign _GEN_394 = 9'h189 == cnt[8:0] ? $signed(-32'shbebc) : $signed(_GEN_393); // @[FFT.scala 34:12]
  assign _GEN_395 = 9'h18a == cnt[8:0] ? $signed(-32'shbfc7) : $signed(_GEN_394); // @[FFT.scala 34:12]
  assign _GEN_396 = 9'h18b == cnt[8:0] ? $signed(-32'shc0d1) : $signed(_GEN_395); // @[FFT.scala 34:12]
  assign _GEN_397 = 9'h18c == cnt[8:0] ? $signed(-32'shc1d8) : $signed(_GEN_396); // @[FFT.scala 34:12]
  assign _GEN_398 = 9'h18d == cnt[8:0] ? $signed(-32'shc2de) : $signed(_GEN_397); // @[FFT.scala 34:12]
  assign _GEN_399 = 9'h18e == cnt[8:0] ? $signed(-32'shc3e2) : $signed(_GEN_398); // @[FFT.scala 34:12]
  assign _GEN_400 = 9'h18f == cnt[8:0] ? $signed(-32'shc4e4) : $signed(_GEN_399); // @[FFT.scala 34:12]
  assign _GEN_401 = 9'h190 == cnt[8:0] ? $signed(-32'shc5e4) : $signed(_GEN_400); // @[FFT.scala 34:12]
  assign _GEN_402 = 9'h191 == cnt[8:0] ? $signed(-32'shc6e2) : $signed(_GEN_401); // @[FFT.scala 34:12]
  assign _GEN_403 = 9'h192 == cnt[8:0] ? $signed(-32'shc7de) : $signed(_GEN_402); // @[FFT.scala 34:12]
  assign _GEN_404 = 9'h193 == cnt[8:0] ? $signed(-32'shc8d9) : $signed(_GEN_403); // @[FFT.scala 34:12]
  assign _GEN_405 = 9'h194 == cnt[8:0] ? $signed(-32'shc9d1) : $signed(_GEN_404); // @[FFT.scala 34:12]
  assign _GEN_406 = 9'h195 == cnt[8:0] ? $signed(-32'shcac7) : $signed(_GEN_405); // @[FFT.scala 34:12]
  assign _GEN_407 = 9'h196 == cnt[8:0] ? $signed(-32'shcbbc) : $signed(_GEN_406); // @[FFT.scala 34:12]
  assign _GEN_408 = 9'h197 == cnt[8:0] ? $signed(-32'shccae) : $signed(_GEN_407); // @[FFT.scala 34:12]
  assign _GEN_409 = 9'h198 == cnt[8:0] ? $signed(-32'shcd9f) : $signed(_GEN_408); // @[FFT.scala 34:12]
  assign _GEN_410 = 9'h199 == cnt[8:0] ? $signed(-32'shce8e) : $signed(_GEN_409); // @[FFT.scala 34:12]
  assign _GEN_411 = 9'h19a == cnt[8:0] ? $signed(-32'shcf7a) : $signed(_GEN_410); // @[FFT.scala 34:12]
  assign _GEN_412 = 9'h19b == cnt[8:0] ? $signed(-32'shd065) : $signed(_GEN_411); // @[FFT.scala 34:12]
  assign _GEN_413 = 9'h19c == cnt[8:0] ? $signed(-32'shd14d) : $signed(_GEN_412); // @[FFT.scala 34:12]
  assign _GEN_414 = 9'h19d == cnt[8:0] ? $signed(-32'shd234) : $signed(_GEN_413); // @[FFT.scala 34:12]
  assign _GEN_415 = 9'h19e == cnt[8:0] ? $signed(-32'shd318) : $signed(_GEN_414); // @[FFT.scala 34:12]
  assign _GEN_416 = 9'h19f == cnt[8:0] ? $signed(-32'shd3fb) : $signed(_GEN_415); // @[FFT.scala 34:12]
  assign _GEN_417 = 9'h1a0 == cnt[8:0] ? $signed(-32'shd4db) : $signed(_GEN_416); // @[FFT.scala 34:12]
  assign _GEN_418 = 9'h1a1 == cnt[8:0] ? $signed(-32'shd5ba) : $signed(_GEN_417); // @[FFT.scala 34:12]
  assign _GEN_419 = 9'h1a2 == cnt[8:0] ? $signed(-32'shd696) : $signed(_GEN_418); // @[FFT.scala 34:12]
  assign _GEN_420 = 9'h1a3 == cnt[8:0] ? $signed(-32'shd770) : $signed(_GEN_419); // @[FFT.scala 34:12]
  assign _GEN_421 = 9'h1a4 == cnt[8:0] ? $signed(-32'shd848) : $signed(_GEN_420); // @[FFT.scala 34:12]
  assign _GEN_422 = 9'h1a5 == cnt[8:0] ? $signed(-32'shd91e) : $signed(_GEN_421); // @[FFT.scala 34:12]
  assign _GEN_423 = 9'h1a6 == cnt[8:0] ? $signed(-32'shd9f2) : $signed(_GEN_422); // @[FFT.scala 34:12]
  assign _GEN_424 = 9'h1a7 == cnt[8:0] ? $signed(-32'shdac4) : $signed(_GEN_423); // @[FFT.scala 34:12]
  assign _GEN_425 = 9'h1a8 == cnt[8:0] ? $signed(-32'shdb94) : $signed(_GEN_424); // @[FFT.scala 34:12]
  assign _GEN_426 = 9'h1a9 == cnt[8:0] ? $signed(-32'shdc62) : $signed(_GEN_425); // @[FFT.scala 34:12]
  assign _GEN_427 = 9'h1aa == cnt[8:0] ? $signed(-32'shdd2d) : $signed(_GEN_426); // @[FFT.scala 34:12]
  assign _GEN_428 = 9'h1ab == cnt[8:0] ? $signed(-32'shddf7) : $signed(_GEN_427); // @[FFT.scala 34:12]
  assign _GEN_429 = 9'h1ac == cnt[8:0] ? $signed(-32'shdebe) : $signed(_GEN_428); // @[FFT.scala 34:12]
  assign _GEN_430 = 9'h1ad == cnt[8:0] ? $signed(-32'shdf83) : $signed(_GEN_429); // @[FFT.scala 34:12]
  assign _GEN_431 = 9'h1ae == cnt[8:0] ? $signed(-32'she046) : $signed(_GEN_430); // @[FFT.scala 34:12]
  assign _GEN_432 = 9'h1af == cnt[8:0] ? $signed(-32'she107) : $signed(_GEN_431); // @[FFT.scala 34:12]
  assign _GEN_433 = 9'h1b0 == cnt[8:0] ? $signed(-32'she1c6) : $signed(_GEN_432); // @[FFT.scala 34:12]
  assign _GEN_434 = 9'h1b1 == cnt[8:0] ? $signed(-32'she282) : $signed(_GEN_433); // @[FFT.scala 34:12]
  assign _GEN_435 = 9'h1b2 == cnt[8:0] ? $signed(-32'she33c) : $signed(_GEN_434); // @[FFT.scala 34:12]
  assign _GEN_436 = 9'h1b3 == cnt[8:0] ? $signed(-32'she3f4) : $signed(_GEN_435); // @[FFT.scala 34:12]
  assign _GEN_437 = 9'h1b4 == cnt[8:0] ? $signed(-32'she4aa) : $signed(_GEN_436); // @[FFT.scala 34:12]
  assign _GEN_438 = 9'h1b5 == cnt[8:0] ? $signed(-32'she55e) : $signed(_GEN_437); // @[FFT.scala 34:12]
  assign _GEN_439 = 9'h1b6 == cnt[8:0] ? $signed(-32'she610) : $signed(_GEN_438); // @[FFT.scala 34:12]
  assign _GEN_440 = 9'h1b7 == cnt[8:0] ? $signed(-32'she6bf) : $signed(_GEN_439); // @[FFT.scala 34:12]
  assign _GEN_441 = 9'h1b8 == cnt[8:0] ? $signed(-32'she76c) : $signed(_GEN_440); // @[FFT.scala 34:12]
  assign _GEN_442 = 9'h1b9 == cnt[8:0] ? $signed(-32'she817) : $signed(_GEN_441); // @[FFT.scala 34:12]
  assign _GEN_443 = 9'h1ba == cnt[8:0] ? $signed(-32'she8bf) : $signed(_GEN_442); // @[FFT.scala 34:12]
  assign _GEN_444 = 9'h1bb == cnt[8:0] ? $signed(-32'she966) : $signed(_GEN_443); // @[FFT.scala 34:12]
  assign _GEN_445 = 9'h1bc == cnt[8:0] ? $signed(-32'shea0a) : $signed(_GEN_444); // @[FFT.scala 34:12]
  assign _GEN_446 = 9'h1bd == cnt[8:0] ? $signed(-32'sheaab) : $signed(_GEN_445); // @[FFT.scala 34:12]
  assign _GEN_447 = 9'h1be == cnt[8:0] ? $signed(-32'sheb4b) : $signed(_GEN_446); // @[FFT.scala 34:12]
  assign _GEN_448 = 9'h1bf == cnt[8:0] ? $signed(-32'shebe8) : $signed(_GEN_447); // @[FFT.scala 34:12]
  assign _GEN_449 = 9'h1c0 == cnt[8:0] ? $signed(-32'shec83) : $signed(_GEN_448); // @[FFT.scala 34:12]
  assign _GEN_450 = 9'h1c1 == cnt[8:0] ? $signed(-32'shed1c) : $signed(_GEN_449); // @[FFT.scala 34:12]
  assign _GEN_451 = 9'h1c2 == cnt[8:0] ? $signed(-32'shedb3) : $signed(_GEN_450); // @[FFT.scala 34:12]
  assign _GEN_452 = 9'h1c3 == cnt[8:0] ? $signed(-32'shee47) : $signed(_GEN_451); // @[FFT.scala 34:12]
  assign _GEN_453 = 9'h1c4 == cnt[8:0] ? $signed(-32'sheed9) : $signed(_GEN_452); // @[FFT.scala 34:12]
  assign _GEN_454 = 9'h1c5 == cnt[8:0] ? $signed(-32'shef68) : $signed(_GEN_453); // @[FFT.scala 34:12]
  assign _GEN_455 = 9'h1c6 == cnt[8:0] ? $signed(-32'sheff5) : $signed(_GEN_454); // @[FFT.scala 34:12]
  assign _GEN_456 = 9'h1c7 == cnt[8:0] ? $signed(-32'shf080) : $signed(_GEN_455); // @[FFT.scala 34:12]
  assign _GEN_457 = 9'h1c8 == cnt[8:0] ? $signed(-32'shf109) : $signed(_GEN_456); // @[FFT.scala 34:12]
  assign _GEN_458 = 9'h1c9 == cnt[8:0] ? $signed(-32'shf18f) : $signed(_GEN_457); // @[FFT.scala 34:12]
  assign _GEN_459 = 9'h1ca == cnt[8:0] ? $signed(-32'shf213) : $signed(_GEN_458); // @[FFT.scala 34:12]
  assign _GEN_460 = 9'h1cb == cnt[8:0] ? $signed(-32'shf295) : $signed(_GEN_459); // @[FFT.scala 34:12]
  assign _GEN_461 = 9'h1cc == cnt[8:0] ? $signed(-32'shf314) : $signed(_GEN_460); // @[FFT.scala 34:12]
  assign _GEN_462 = 9'h1cd == cnt[8:0] ? $signed(-32'shf391) : $signed(_GEN_461); // @[FFT.scala 34:12]
  assign _GEN_463 = 9'h1ce == cnt[8:0] ? $signed(-32'shf40c) : $signed(_GEN_462); // @[FFT.scala 34:12]
  assign _GEN_464 = 9'h1cf == cnt[8:0] ? $signed(-32'shf484) : $signed(_GEN_463); // @[FFT.scala 34:12]
  assign _GEN_465 = 9'h1d0 == cnt[8:0] ? $signed(-32'shf4fa) : $signed(_GEN_464); // @[FFT.scala 34:12]
  assign _GEN_466 = 9'h1d1 == cnt[8:0] ? $signed(-32'shf56e) : $signed(_GEN_465); // @[FFT.scala 34:12]
  assign _GEN_467 = 9'h1d2 == cnt[8:0] ? $signed(-32'shf5df) : $signed(_GEN_466); // @[FFT.scala 34:12]
  assign _GEN_468 = 9'h1d3 == cnt[8:0] ? $signed(-32'shf64e) : $signed(_GEN_467); // @[FFT.scala 34:12]
  assign _GEN_469 = 9'h1d4 == cnt[8:0] ? $signed(-32'shf6ba) : $signed(_GEN_468); // @[FFT.scala 34:12]
  assign _GEN_470 = 9'h1d5 == cnt[8:0] ? $signed(-32'shf724) : $signed(_GEN_469); // @[FFT.scala 34:12]
  assign _GEN_471 = 9'h1d6 == cnt[8:0] ? $signed(-32'shf78c) : $signed(_GEN_470); // @[FFT.scala 34:12]
  assign _GEN_472 = 9'h1d7 == cnt[8:0] ? $signed(-32'shf7f1) : $signed(_GEN_471); // @[FFT.scala 34:12]
  assign _GEN_473 = 9'h1d8 == cnt[8:0] ? $signed(-32'shf854) : $signed(_GEN_472); // @[FFT.scala 34:12]
  assign _GEN_474 = 9'h1d9 == cnt[8:0] ? $signed(-32'shf8b4) : $signed(_GEN_473); // @[FFT.scala 34:12]
  assign _GEN_475 = 9'h1da == cnt[8:0] ? $signed(-32'shf913) : $signed(_GEN_474); // @[FFT.scala 34:12]
  assign _GEN_476 = 9'h1db == cnt[8:0] ? $signed(-32'shf96e) : $signed(_GEN_475); // @[FFT.scala 34:12]
  assign _GEN_477 = 9'h1dc == cnt[8:0] ? $signed(-32'shf9c8) : $signed(_GEN_476); // @[FFT.scala 34:12]
  assign _GEN_478 = 9'h1dd == cnt[8:0] ? $signed(-32'shfa1f) : $signed(_GEN_477); // @[FFT.scala 34:12]
  assign _GEN_479 = 9'h1de == cnt[8:0] ? $signed(-32'shfa73) : $signed(_GEN_478); // @[FFT.scala 34:12]
  assign _GEN_480 = 9'h1df == cnt[8:0] ? $signed(-32'shfac5) : $signed(_GEN_479); // @[FFT.scala 34:12]
  assign _GEN_481 = 9'h1e0 == cnt[8:0] ? $signed(-32'shfb15) : $signed(_GEN_480); // @[FFT.scala 34:12]
  assign _GEN_482 = 9'h1e1 == cnt[8:0] ? $signed(-32'shfb62) : $signed(_GEN_481); // @[FFT.scala 34:12]
  assign _GEN_483 = 9'h1e2 == cnt[8:0] ? $signed(-32'shfbad) : $signed(_GEN_482); // @[FFT.scala 34:12]
  assign _GEN_484 = 9'h1e3 == cnt[8:0] ? $signed(-32'shfbf5) : $signed(_GEN_483); // @[FFT.scala 34:12]
  assign _GEN_485 = 9'h1e4 == cnt[8:0] ? $signed(-32'shfc3b) : $signed(_GEN_484); // @[FFT.scala 34:12]
  assign _GEN_486 = 9'h1e5 == cnt[8:0] ? $signed(-32'shfc7f) : $signed(_GEN_485); // @[FFT.scala 34:12]
  assign _GEN_487 = 9'h1e6 == cnt[8:0] ? $signed(-32'shfcc0) : $signed(_GEN_486); // @[FFT.scala 34:12]
  assign _GEN_488 = 9'h1e7 == cnt[8:0] ? $signed(-32'shfcfe) : $signed(_GEN_487); // @[FFT.scala 34:12]
  assign _GEN_489 = 9'h1e8 == cnt[8:0] ? $signed(-32'shfd3b) : $signed(_GEN_488); // @[FFT.scala 34:12]
  assign _GEN_490 = 9'h1e9 == cnt[8:0] ? $signed(-32'shfd74) : $signed(_GEN_489); // @[FFT.scala 34:12]
  assign _GEN_491 = 9'h1ea == cnt[8:0] ? $signed(-32'shfdac) : $signed(_GEN_490); // @[FFT.scala 34:12]
  assign _GEN_492 = 9'h1eb == cnt[8:0] ? $signed(-32'shfde1) : $signed(_GEN_491); // @[FFT.scala 34:12]
  assign _GEN_493 = 9'h1ec == cnt[8:0] ? $signed(-32'shfe13) : $signed(_GEN_492); // @[FFT.scala 34:12]
  assign _GEN_494 = 9'h1ed == cnt[8:0] ? $signed(-32'shfe43) : $signed(_GEN_493); // @[FFT.scala 34:12]
  assign _GEN_495 = 9'h1ee == cnt[8:0] ? $signed(-32'shfe71) : $signed(_GEN_494); // @[FFT.scala 34:12]
  assign _GEN_496 = 9'h1ef == cnt[8:0] ? $signed(-32'shfe9c) : $signed(_GEN_495); // @[FFT.scala 34:12]
  assign _GEN_497 = 9'h1f0 == cnt[8:0] ? $signed(-32'shfec4) : $signed(_GEN_496); // @[FFT.scala 34:12]
  assign _GEN_498 = 9'h1f1 == cnt[8:0] ? $signed(-32'shfeeb) : $signed(_GEN_497); // @[FFT.scala 34:12]
  assign _GEN_499 = 9'h1f2 == cnt[8:0] ? $signed(-32'shff0e) : $signed(_GEN_498); // @[FFT.scala 34:12]
  assign _GEN_500 = 9'h1f3 == cnt[8:0] ? $signed(-32'shff30) : $signed(_GEN_499); // @[FFT.scala 34:12]
  assign _GEN_501 = 9'h1f4 == cnt[8:0] ? $signed(-32'shff4e) : $signed(_GEN_500); // @[FFT.scala 34:12]
  assign _GEN_502 = 9'h1f5 == cnt[8:0] ? $signed(-32'shff6b) : $signed(_GEN_501); // @[FFT.scala 34:12]
  assign _GEN_503 = 9'h1f6 == cnt[8:0] ? $signed(-32'shff85) : $signed(_GEN_502); // @[FFT.scala 34:12]
  assign _GEN_504 = 9'h1f7 == cnt[8:0] ? $signed(-32'shff9c) : $signed(_GEN_503); // @[FFT.scala 34:12]
  assign _GEN_505 = 9'h1f8 == cnt[8:0] ? $signed(-32'shffb1) : $signed(_GEN_504); // @[FFT.scala 34:12]
  assign _GEN_506 = 9'h1f9 == cnt[8:0] ? $signed(-32'shffc4) : $signed(_GEN_505); // @[FFT.scala 34:12]
  assign _GEN_507 = 9'h1fa == cnt[8:0] ? $signed(-32'shffd4) : $signed(_GEN_506); // @[FFT.scala 34:12]
  assign _GEN_508 = 9'h1fb == cnt[8:0] ? $signed(-32'shffe1) : $signed(_GEN_507); // @[FFT.scala 34:12]
  assign _GEN_509 = 9'h1fc == cnt[8:0] ? $signed(-32'shffec) : $signed(_GEN_508); // @[FFT.scala 34:12]
  assign _GEN_510 = 9'h1fd == cnt[8:0] ? $signed(-32'shfff5) : $signed(_GEN_509); // @[FFT.scala 34:12]
  assign _GEN_511 = 9'h1fe == cnt[8:0] ? $signed(-32'shfffb) : $signed(_GEN_510); // @[FFT.scala 34:12]
  assign _GEN_514 = 9'h1 == cnt[8:0] ? $signed(-32'sh192) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_515 = 9'h2 == cnt[8:0] ? $signed(-32'sh324) : $signed(_GEN_514); // @[FFT.scala 35:12]
  assign _GEN_516 = 9'h3 == cnt[8:0] ? $signed(-32'sh4b6) : $signed(_GEN_515); // @[FFT.scala 35:12]
  assign _GEN_517 = 9'h4 == cnt[8:0] ? $signed(-32'sh648) : $signed(_GEN_516); // @[FFT.scala 35:12]
  assign _GEN_518 = 9'h5 == cnt[8:0] ? $signed(-32'sh7da) : $signed(_GEN_517); // @[FFT.scala 35:12]
  assign _GEN_519 = 9'h6 == cnt[8:0] ? $signed(-32'sh96c) : $signed(_GEN_518); // @[FFT.scala 35:12]
  assign _GEN_520 = 9'h7 == cnt[8:0] ? $signed(-32'shafe) : $signed(_GEN_519); // @[FFT.scala 35:12]
  assign _GEN_521 = 9'h8 == cnt[8:0] ? $signed(-32'shc90) : $signed(_GEN_520); // @[FFT.scala 35:12]
  assign _GEN_522 = 9'h9 == cnt[8:0] ? $signed(-32'she21) : $signed(_GEN_521); // @[FFT.scala 35:12]
  assign _GEN_523 = 9'ha == cnt[8:0] ? $signed(-32'shfb3) : $signed(_GEN_522); // @[FFT.scala 35:12]
  assign _GEN_524 = 9'hb == cnt[8:0] ? $signed(-32'sh1144) : $signed(_GEN_523); // @[FFT.scala 35:12]
  assign _GEN_525 = 9'hc == cnt[8:0] ? $signed(-32'sh12d5) : $signed(_GEN_524); // @[FFT.scala 35:12]
  assign _GEN_526 = 9'hd == cnt[8:0] ? $signed(-32'sh1466) : $signed(_GEN_525); // @[FFT.scala 35:12]
  assign _GEN_527 = 9'he == cnt[8:0] ? $signed(-32'sh15f7) : $signed(_GEN_526); // @[FFT.scala 35:12]
  assign _GEN_528 = 9'hf == cnt[8:0] ? $signed(-32'sh1787) : $signed(_GEN_527); // @[FFT.scala 35:12]
  assign _GEN_529 = 9'h10 == cnt[8:0] ? $signed(-32'sh1918) : $signed(_GEN_528); // @[FFT.scala 35:12]
  assign _GEN_530 = 9'h11 == cnt[8:0] ? $signed(-32'sh1aa8) : $signed(_GEN_529); // @[FFT.scala 35:12]
  assign _GEN_531 = 9'h12 == cnt[8:0] ? $signed(-32'sh1c38) : $signed(_GEN_530); // @[FFT.scala 35:12]
  assign _GEN_532 = 9'h13 == cnt[8:0] ? $signed(-32'sh1dc7) : $signed(_GEN_531); // @[FFT.scala 35:12]
  assign _GEN_533 = 9'h14 == cnt[8:0] ? $signed(-32'sh1f56) : $signed(_GEN_532); // @[FFT.scala 35:12]
  assign _GEN_534 = 9'h15 == cnt[8:0] ? $signed(-32'sh20e5) : $signed(_GEN_533); // @[FFT.scala 35:12]
  assign _GEN_535 = 9'h16 == cnt[8:0] ? $signed(-32'sh2274) : $signed(_GEN_534); // @[FFT.scala 35:12]
  assign _GEN_536 = 9'h17 == cnt[8:0] ? $signed(-32'sh2402) : $signed(_GEN_535); // @[FFT.scala 35:12]
  assign _GEN_537 = 9'h18 == cnt[8:0] ? $signed(-32'sh2590) : $signed(_GEN_536); // @[FFT.scala 35:12]
  assign _GEN_538 = 9'h19 == cnt[8:0] ? $signed(-32'sh271e) : $signed(_GEN_537); // @[FFT.scala 35:12]
  assign _GEN_539 = 9'h1a == cnt[8:0] ? $signed(-32'sh28ab) : $signed(_GEN_538); // @[FFT.scala 35:12]
  assign _GEN_540 = 9'h1b == cnt[8:0] ? $signed(-32'sh2a38) : $signed(_GEN_539); // @[FFT.scala 35:12]
  assign _GEN_541 = 9'h1c == cnt[8:0] ? $signed(-32'sh2bc4) : $signed(_GEN_540); // @[FFT.scala 35:12]
  assign _GEN_542 = 9'h1d == cnt[8:0] ? $signed(-32'sh2d50) : $signed(_GEN_541); // @[FFT.scala 35:12]
  assign _GEN_543 = 9'h1e == cnt[8:0] ? $signed(-32'sh2edc) : $signed(_GEN_542); // @[FFT.scala 35:12]
  assign _GEN_544 = 9'h1f == cnt[8:0] ? $signed(-32'sh3067) : $signed(_GEN_543); // @[FFT.scala 35:12]
  assign _GEN_545 = 9'h20 == cnt[8:0] ? $signed(-32'sh31f1) : $signed(_GEN_544); // @[FFT.scala 35:12]
  assign _GEN_546 = 9'h21 == cnt[8:0] ? $signed(-32'sh337c) : $signed(_GEN_545); // @[FFT.scala 35:12]
  assign _GEN_547 = 9'h22 == cnt[8:0] ? $signed(-32'sh3505) : $signed(_GEN_546); // @[FFT.scala 35:12]
  assign _GEN_548 = 9'h23 == cnt[8:0] ? $signed(-32'sh368e) : $signed(_GEN_547); // @[FFT.scala 35:12]
  assign _GEN_549 = 9'h24 == cnt[8:0] ? $signed(-32'sh3817) : $signed(_GEN_548); // @[FFT.scala 35:12]
  assign _GEN_550 = 9'h25 == cnt[8:0] ? $signed(-32'sh399f) : $signed(_GEN_549); // @[FFT.scala 35:12]
  assign _GEN_551 = 9'h26 == cnt[8:0] ? $signed(-32'sh3b27) : $signed(_GEN_550); // @[FFT.scala 35:12]
  assign _GEN_552 = 9'h27 == cnt[8:0] ? $signed(-32'sh3cae) : $signed(_GEN_551); // @[FFT.scala 35:12]
  assign _GEN_553 = 9'h28 == cnt[8:0] ? $signed(-32'sh3e34) : $signed(_GEN_552); // @[FFT.scala 35:12]
  assign _GEN_554 = 9'h29 == cnt[8:0] ? $signed(-32'sh3fba) : $signed(_GEN_553); // @[FFT.scala 35:12]
  assign _GEN_555 = 9'h2a == cnt[8:0] ? $signed(-32'sh413f) : $signed(_GEN_554); // @[FFT.scala 35:12]
  assign _GEN_556 = 9'h2b == cnt[8:0] ? $signed(-32'sh42c3) : $signed(_GEN_555); // @[FFT.scala 35:12]
  assign _GEN_557 = 9'h2c == cnt[8:0] ? $signed(-32'sh4447) : $signed(_GEN_556); // @[FFT.scala 35:12]
  assign _GEN_558 = 9'h2d == cnt[8:0] ? $signed(-32'sh45cb) : $signed(_GEN_557); // @[FFT.scala 35:12]
  assign _GEN_559 = 9'h2e == cnt[8:0] ? $signed(-32'sh474d) : $signed(_GEN_558); // @[FFT.scala 35:12]
  assign _GEN_560 = 9'h2f == cnt[8:0] ? $signed(-32'sh48cf) : $signed(_GEN_559); // @[FFT.scala 35:12]
  assign _GEN_561 = 9'h30 == cnt[8:0] ? $signed(-32'sh4a50) : $signed(_GEN_560); // @[FFT.scala 35:12]
  assign _GEN_562 = 9'h31 == cnt[8:0] ? $signed(-32'sh4bd1) : $signed(_GEN_561); // @[FFT.scala 35:12]
  assign _GEN_563 = 9'h32 == cnt[8:0] ? $signed(-32'sh4d50) : $signed(_GEN_562); // @[FFT.scala 35:12]
  assign _GEN_564 = 9'h33 == cnt[8:0] ? $signed(-32'sh4ecf) : $signed(_GEN_563); // @[FFT.scala 35:12]
  assign _GEN_565 = 9'h34 == cnt[8:0] ? $signed(-32'sh504d) : $signed(_GEN_564); // @[FFT.scala 35:12]
  assign _GEN_566 = 9'h35 == cnt[8:0] ? $signed(-32'sh51cb) : $signed(_GEN_565); // @[FFT.scala 35:12]
  assign _GEN_567 = 9'h36 == cnt[8:0] ? $signed(-32'sh5348) : $signed(_GEN_566); // @[FFT.scala 35:12]
  assign _GEN_568 = 9'h37 == cnt[8:0] ? $signed(-32'sh54c3) : $signed(_GEN_567); // @[FFT.scala 35:12]
  assign _GEN_569 = 9'h38 == cnt[8:0] ? $signed(-32'sh563e) : $signed(_GEN_568); // @[FFT.scala 35:12]
  assign _GEN_570 = 9'h39 == cnt[8:0] ? $signed(-32'sh57b9) : $signed(_GEN_569); // @[FFT.scala 35:12]
  assign _GEN_571 = 9'h3a == cnt[8:0] ? $signed(-32'sh5932) : $signed(_GEN_570); // @[FFT.scala 35:12]
  assign _GEN_572 = 9'h3b == cnt[8:0] ? $signed(-32'sh5aaa) : $signed(_GEN_571); // @[FFT.scala 35:12]
  assign _GEN_573 = 9'h3c == cnt[8:0] ? $signed(-32'sh5c22) : $signed(_GEN_572); // @[FFT.scala 35:12]
  assign _GEN_574 = 9'h3d == cnt[8:0] ? $signed(-32'sh5d99) : $signed(_GEN_573); // @[FFT.scala 35:12]
  assign _GEN_575 = 9'h3e == cnt[8:0] ? $signed(-32'sh5f0f) : $signed(_GEN_574); // @[FFT.scala 35:12]
  assign _GEN_576 = 9'h3f == cnt[8:0] ? $signed(-32'sh6084) : $signed(_GEN_575); // @[FFT.scala 35:12]
  assign _GEN_577 = 9'h40 == cnt[8:0] ? $signed(-32'sh61f8) : $signed(_GEN_576); // @[FFT.scala 35:12]
  assign _GEN_578 = 9'h41 == cnt[8:0] ? $signed(-32'sh636b) : $signed(_GEN_577); // @[FFT.scala 35:12]
  assign _GEN_579 = 9'h42 == cnt[8:0] ? $signed(-32'sh64dd) : $signed(_GEN_578); // @[FFT.scala 35:12]
  assign _GEN_580 = 9'h43 == cnt[8:0] ? $signed(-32'sh664e) : $signed(_GEN_579); // @[FFT.scala 35:12]
  assign _GEN_581 = 9'h44 == cnt[8:0] ? $signed(-32'sh67be) : $signed(_GEN_580); // @[FFT.scala 35:12]
  assign _GEN_582 = 9'h45 == cnt[8:0] ? $signed(-32'sh692d) : $signed(_GEN_581); // @[FFT.scala 35:12]
  assign _GEN_583 = 9'h46 == cnt[8:0] ? $signed(-32'sh6a9b) : $signed(_GEN_582); // @[FFT.scala 35:12]
  assign _GEN_584 = 9'h47 == cnt[8:0] ? $signed(-32'sh6c08) : $signed(_GEN_583); // @[FFT.scala 35:12]
  assign _GEN_585 = 9'h48 == cnt[8:0] ? $signed(-32'sh6d74) : $signed(_GEN_584); // @[FFT.scala 35:12]
  assign _GEN_586 = 9'h49 == cnt[8:0] ? $signed(-32'sh6edf) : $signed(_GEN_585); // @[FFT.scala 35:12]
  assign _GEN_587 = 9'h4a == cnt[8:0] ? $signed(-32'sh7049) : $signed(_GEN_586); // @[FFT.scala 35:12]
  assign _GEN_588 = 9'h4b == cnt[8:0] ? $signed(-32'sh71b2) : $signed(_GEN_587); // @[FFT.scala 35:12]
  assign _GEN_589 = 9'h4c == cnt[8:0] ? $signed(-32'sh731a) : $signed(_GEN_588); // @[FFT.scala 35:12]
  assign _GEN_590 = 9'h4d == cnt[8:0] ? $signed(-32'sh7480) : $signed(_GEN_589); // @[FFT.scala 35:12]
  assign _GEN_591 = 9'h4e == cnt[8:0] ? $signed(-32'sh75e6) : $signed(_GEN_590); // @[FFT.scala 35:12]
  assign _GEN_592 = 9'h4f == cnt[8:0] ? $signed(-32'sh774a) : $signed(_GEN_591); // @[FFT.scala 35:12]
  assign _GEN_593 = 9'h50 == cnt[8:0] ? $signed(-32'sh78ad) : $signed(_GEN_592); // @[FFT.scala 35:12]
  assign _GEN_594 = 9'h51 == cnt[8:0] ? $signed(-32'sh7a10) : $signed(_GEN_593); // @[FFT.scala 35:12]
  assign _GEN_595 = 9'h52 == cnt[8:0] ? $signed(-32'sh7b70) : $signed(_GEN_594); // @[FFT.scala 35:12]
  assign _GEN_596 = 9'h53 == cnt[8:0] ? $signed(-32'sh7cd0) : $signed(_GEN_595); // @[FFT.scala 35:12]
  assign _GEN_597 = 9'h54 == cnt[8:0] ? $signed(-32'sh7e2f) : $signed(_GEN_596); // @[FFT.scala 35:12]
  assign _GEN_598 = 9'h55 == cnt[8:0] ? $signed(-32'sh7f8c) : $signed(_GEN_597); // @[FFT.scala 35:12]
  assign _GEN_599 = 9'h56 == cnt[8:0] ? $signed(-32'sh80e8) : $signed(_GEN_598); // @[FFT.scala 35:12]
  assign _GEN_600 = 9'h57 == cnt[8:0] ? $signed(-32'sh8243) : $signed(_GEN_599); // @[FFT.scala 35:12]
  assign _GEN_601 = 9'h58 == cnt[8:0] ? $signed(-32'sh839c) : $signed(_GEN_600); // @[FFT.scala 35:12]
  assign _GEN_602 = 9'h59 == cnt[8:0] ? $signed(-32'sh84f5) : $signed(_GEN_601); // @[FFT.scala 35:12]
  assign _GEN_603 = 9'h5a == cnt[8:0] ? $signed(-32'sh864c) : $signed(_GEN_602); // @[FFT.scala 35:12]
  assign _GEN_604 = 9'h5b == cnt[8:0] ? $signed(-32'sh87a1) : $signed(_GEN_603); // @[FFT.scala 35:12]
  assign _GEN_605 = 9'h5c == cnt[8:0] ? $signed(-32'sh88f6) : $signed(_GEN_604); // @[FFT.scala 35:12]
  assign _GEN_606 = 9'h5d == cnt[8:0] ? $signed(-32'sh8a49) : $signed(_GEN_605); // @[FFT.scala 35:12]
  assign _GEN_607 = 9'h5e == cnt[8:0] ? $signed(-32'sh8b9a) : $signed(_GEN_606); // @[FFT.scala 35:12]
  assign _GEN_608 = 9'h5f == cnt[8:0] ? $signed(-32'sh8ceb) : $signed(_GEN_607); // @[FFT.scala 35:12]
  assign _GEN_609 = 9'h60 == cnt[8:0] ? $signed(-32'sh8e3a) : $signed(_GEN_608); // @[FFT.scala 35:12]
  assign _GEN_610 = 9'h61 == cnt[8:0] ? $signed(-32'sh8f88) : $signed(_GEN_609); // @[FFT.scala 35:12]
  assign _GEN_611 = 9'h62 == cnt[8:0] ? $signed(-32'sh90d4) : $signed(_GEN_610); // @[FFT.scala 35:12]
  assign _GEN_612 = 9'h63 == cnt[8:0] ? $signed(-32'sh921f) : $signed(_GEN_611); // @[FFT.scala 35:12]
  assign _GEN_613 = 9'h64 == cnt[8:0] ? $signed(-32'sh9368) : $signed(_GEN_612); // @[FFT.scala 35:12]
  assign _GEN_614 = 9'h65 == cnt[8:0] ? $signed(-32'sh94b0) : $signed(_GEN_613); // @[FFT.scala 35:12]
  assign _GEN_615 = 9'h66 == cnt[8:0] ? $signed(-32'sh95f7) : $signed(_GEN_614); // @[FFT.scala 35:12]
  assign _GEN_616 = 9'h67 == cnt[8:0] ? $signed(-32'sh973c) : $signed(_GEN_615); // @[FFT.scala 35:12]
  assign _GEN_617 = 9'h68 == cnt[8:0] ? $signed(-32'sh9880) : $signed(_GEN_616); // @[FFT.scala 35:12]
  assign _GEN_618 = 9'h69 == cnt[8:0] ? $signed(-32'sh99c2) : $signed(_GEN_617); // @[FFT.scala 35:12]
  assign _GEN_619 = 9'h6a == cnt[8:0] ? $signed(-32'sh9b03) : $signed(_GEN_618); // @[FFT.scala 35:12]
  assign _GEN_620 = 9'h6b == cnt[8:0] ? $signed(-32'sh9c42) : $signed(_GEN_619); // @[FFT.scala 35:12]
  assign _GEN_621 = 9'h6c == cnt[8:0] ? $signed(-32'sh9d80) : $signed(_GEN_620); // @[FFT.scala 35:12]
  assign _GEN_622 = 9'h6d == cnt[8:0] ? $signed(-32'sh9ebc) : $signed(_GEN_621); // @[FFT.scala 35:12]
  assign _GEN_623 = 9'h6e == cnt[8:0] ? $signed(-32'sh9ff7) : $signed(_GEN_622); // @[FFT.scala 35:12]
  assign _GEN_624 = 9'h6f == cnt[8:0] ? $signed(-32'sha130) : $signed(_GEN_623); // @[FFT.scala 35:12]
  assign _GEN_625 = 9'h70 == cnt[8:0] ? $signed(-32'sha268) : $signed(_GEN_624); // @[FFT.scala 35:12]
  assign _GEN_626 = 9'h71 == cnt[8:0] ? $signed(-32'sha39e) : $signed(_GEN_625); // @[FFT.scala 35:12]
  assign _GEN_627 = 9'h72 == cnt[8:0] ? $signed(-32'sha4d2) : $signed(_GEN_626); // @[FFT.scala 35:12]
  assign _GEN_628 = 9'h73 == cnt[8:0] ? $signed(-32'sha605) : $signed(_GEN_627); // @[FFT.scala 35:12]
  assign _GEN_629 = 9'h74 == cnt[8:0] ? $signed(-32'sha736) : $signed(_GEN_628); // @[FFT.scala 35:12]
  assign _GEN_630 = 9'h75 == cnt[8:0] ? $signed(-32'sha866) : $signed(_GEN_629); // @[FFT.scala 35:12]
  assign _GEN_631 = 9'h76 == cnt[8:0] ? $signed(-32'sha994) : $signed(_GEN_630); // @[FFT.scala 35:12]
  assign _GEN_632 = 9'h77 == cnt[8:0] ? $signed(-32'shaac1) : $signed(_GEN_631); // @[FFT.scala 35:12]
  assign _GEN_633 = 9'h78 == cnt[8:0] ? $signed(-32'shabeb) : $signed(_GEN_632); // @[FFT.scala 35:12]
  assign _GEN_634 = 9'h79 == cnt[8:0] ? $signed(-32'shad14) : $signed(_GEN_633); // @[FFT.scala 35:12]
  assign _GEN_635 = 9'h7a == cnt[8:0] ? $signed(-32'shae3c) : $signed(_GEN_634); // @[FFT.scala 35:12]
  assign _GEN_636 = 9'h7b == cnt[8:0] ? $signed(-32'shaf62) : $signed(_GEN_635); // @[FFT.scala 35:12]
  assign _GEN_637 = 9'h7c == cnt[8:0] ? $signed(-32'shb086) : $signed(_GEN_636); // @[FFT.scala 35:12]
  assign _GEN_638 = 9'h7d == cnt[8:0] ? $signed(-32'shb1a8) : $signed(_GEN_637); // @[FFT.scala 35:12]
  assign _GEN_639 = 9'h7e == cnt[8:0] ? $signed(-32'shb2c9) : $signed(_GEN_638); // @[FFT.scala 35:12]
  assign _GEN_640 = 9'h7f == cnt[8:0] ? $signed(-32'shb3e8) : $signed(_GEN_639); // @[FFT.scala 35:12]
  assign _GEN_641 = 9'h80 == cnt[8:0] ? $signed(-32'shb505) : $signed(_GEN_640); // @[FFT.scala 35:12]
  assign _GEN_642 = 9'h81 == cnt[8:0] ? $signed(-32'shb620) : $signed(_GEN_641); // @[FFT.scala 35:12]
  assign _GEN_643 = 9'h82 == cnt[8:0] ? $signed(-32'shb73a) : $signed(_GEN_642); // @[FFT.scala 35:12]
  assign _GEN_644 = 9'h83 == cnt[8:0] ? $signed(-32'shb852) : $signed(_GEN_643); // @[FFT.scala 35:12]
  assign _GEN_645 = 9'h84 == cnt[8:0] ? $signed(-32'shb968) : $signed(_GEN_644); // @[FFT.scala 35:12]
  assign _GEN_646 = 9'h85 == cnt[8:0] ? $signed(-32'shba7d) : $signed(_GEN_645); // @[FFT.scala 35:12]
  assign _GEN_647 = 9'h86 == cnt[8:0] ? $signed(-32'shbb8f) : $signed(_GEN_646); // @[FFT.scala 35:12]
  assign _GEN_648 = 9'h87 == cnt[8:0] ? $signed(-32'shbca0) : $signed(_GEN_647); // @[FFT.scala 35:12]
  assign _GEN_649 = 9'h88 == cnt[8:0] ? $signed(-32'shbdaf) : $signed(_GEN_648); // @[FFT.scala 35:12]
  assign _GEN_650 = 9'h89 == cnt[8:0] ? $signed(-32'shbebc) : $signed(_GEN_649); // @[FFT.scala 35:12]
  assign _GEN_651 = 9'h8a == cnt[8:0] ? $signed(-32'shbfc7) : $signed(_GEN_650); // @[FFT.scala 35:12]
  assign _GEN_652 = 9'h8b == cnt[8:0] ? $signed(-32'shc0d1) : $signed(_GEN_651); // @[FFT.scala 35:12]
  assign _GEN_653 = 9'h8c == cnt[8:0] ? $signed(-32'shc1d8) : $signed(_GEN_652); // @[FFT.scala 35:12]
  assign _GEN_654 = 9'h8d == cnt[8:0] ? $signed(-32'shc2de) : $signed(_GEN_653); // @[FFT.scala 35:12]
  assign _GEN_655 = 9'h8e == cnt[8:0] ? $signed(-32'shc3e2) : $signed(_GEN_654); // @[FFT.scala 35:12]
  assign _GEN_656 = 9'h8f == cnt[8:0] ? $signed(-32'shc4e4) : $signed(_GEN_655); // @[FFT.scala 35:12]
  assign _GEN_657 = 9'h90 == cnt[8:0] ? $signed(-32'shc5e4) : $signed(_GEN_656); // @[FFT.scala 35:12]
  assign _GEN_658 = 9'h91 == cnt[8:0] ? $signed(-32'shc6e2) : $signed(_GEN_657); // @[FFT.scala 35:12]
  assign _GEN_659 = 9'h92 == cnt[8:0] ? $signed(-32'shc7de) : $signed(_GEN_658); // @[FFT.scala 35:12]
  assign _GEN_660 = 9'h93 == cnt[8:0] ? $signed(-32'shc8d9) : $signed(_GEN_659); // @[FFT.scala 35:12]
  assign _GEN_661 = 9'h94 == cnt[8:0] ? $signed(-32'shc9d1) : $signed(_GEN_660); // @[FFT.scala 35:12]
  assign _GEN_662 = 9'h95 == cnt[8:0] ? $signed(-32'shcac7) : $signed(_GEN_661); // @[FFT.scala 35:12]
  assign _GEN_663 = 9'h96 == cnt[8:0] ? $signed(-32'shcbbc) : $signed(_GEN_662); // @[FFT.scala 35:12]
  assign _GEN_664 = 9'h97 == cnt[8:0] ? $signed(-32'shccae) : $signed(_GEN_663); // @[FFT.scala 35:12]
  assign _GEN_665 = 9'h98 == cnt[8:0] ? $signed(-32'shcd9f) : $signed(_GEN_664); // @[FFT.scala 35:12]
  assign _GEN_666 = 9'h99 == cnt[8:0] ? $signed(-32'shce8e) : $signed(_GEN_665); // @[FFT.scala 35:12]
  assign _GEN_667 = 9'h9a == cnt[8:0] ? $signed(-32'shcf7a) : $signed(_GEN_666); // @[FFT.scala 35:12]
  assign _GEN_668 = 9'h9b == cnt[8:0] ? $signed(-32'shd065) : $signed(_GEN_667); // @[FFT.scala 35:12]
  assign _GEN_669 = 9'h9c == cnt[8:0] ? $signed(-32'shd14d) : $signed(_GEN_668); // @[FFT.scala 35:12]
  assign _GEN_670 = 9'h9d == cnt[8:0] ? $signed(-32'shd234) : $signed(_GEN_669); // @[FFT.scala 35:12]
  assign _GEN_671 = 9'h9e == cnt[8:0] ? $signed(-32'shd318) : $signed(_GEN_670); // @[FFT.scala 35:12]
  assign _GEN_672 = 9'h9f == cnt[8:0] ? $signed(-32'shd3fb) : $signed(_GEN_671); // @[FFT.scala 35:12]
  assign _GEN_673 = 9'ha0 == cnt[8:0] ? $signed(-32'shd4db) : $signed(_GEN_672); // @[FFT.scala 35:12]
  assign _GEN_674 = 9'ha1 == cnt[8:0] ? $signed(-32'shd5ba) : $signed(_GEN_673); // @[FFT.scala 35:12]
  assign _GEN_675 = 9'ha2 == cnt[8:0] ? $signed(-32'shd696) : $signed(_GEN_674); // @[FFT.scala 35:12]
  assign _GEN_676 = 9'ha3 == cnt[8:0] ? $signed(-32'shd770) : $signed(_GEN_675); // @[FFT.scala 35:12]
  assign _GEN_677 = 9'ha4 == cnt[8:0] ? $signed(-32'shd848) : $signed(_GEN_676); // @[FFT.scala 35:12]
  assign _GEN_678 = 9'ha5 == cnt[8:0] ? $signed(-32'shd91e) : $signed(_GEN_677); // @[FFT.scala 35:12]
  assign _GEN_679 = 9'ha6 == cnt[8:0] ? $signed(-32'shd9f2) : $signed(_GEN_678); // @[FFT.scala 35:12]
  assign _GEN_680 = 9'ha7 == cnt[8:0] ? $signed(-32'shdac4) : $signed(_GEN_679); // @[FFT.scala 35:12]
  assign _GEN_681 = 9'ha8 == cnt[8:0] ? $signed(-32'shdb94) : $signed(_GEN_680); // @[FFT.scala 35:12]
  assign _GEN_682 = 9'ha9 == cnt[8:0] ? $signed(-32'shdc62) : $signed(_GEN_681); // @[FFT.scala 35:12]
  assign _GEN_683 = 9'haa == cnt[8:0] ? $signed(-32'shdd2d) : $signed(_GEN_682); // @[FFT.scala 35:12]
  assign _GEN_684 = 9'hab == cnt[8:0] ? $signed(-32'shddf7) : $signed(_GEN_683); // @[FFT.scala 35:12]
  assign _GEN_685 = 9'hac == cnt[8:0] ? $signed(-32'shdebe) : $signed(_GEN_684); // @[FFT.scala 35:12]
  assign _GEN_686 = 9'had == cnt[8:0] ? $signed(-32'shdf83) : $signed(_GEN_685); // @[FFT.scala 35:12]
  assign _GEN_687 = 9'hae == cnt[8:0] ? $signed(-32'she046) : $signed(_GEN_686); // @[FFT.scala 35:12]
  assign _GEN_688 = 9'haf == cnt[8:0] ? $signed(-32'she107) : $signed(_GEN_687); // @[FFT.scala 35:12]
  assign _GEN_689 = 9'hb0 == cnt[8:0] ? $signed(-32'she1c6) : $signed(_GEN_688); // @[FFT.scala 35:12]
  assign _GEN_690 = 9'hb1 == cnt[8:0] ? $signed(-32'she282) : $signed(_GEN_689); // @[FFT.scala 35:12]
  assign _GEN_691 = 9'hb2 == cnt[8:0] ? $signed(-32'she33c) : $signed(_GEN_690); // @[FFT.scala 35:12]
  assign _GEN_692 = 9'hb3 == cnt[8:0] ? $signed(-32'she3f4) : $signed(_GEN_691); // @[FFT.scala 35:12]
  assign _GEN_693 = 9'hb4 == cnt[8:0] ? $signed(-32'she4aa) : $signed(_GEN_692); // @[FFT.scala 35:12]
  assign _GEN_694 = 9'hb5 == cnt[8:0] ? $signed(-32'she55e) : $signed(_GEN_693); // @[FFT.scala 35:12]
  assign _GEN_695 = 9'hb6 == cnt[8:0] ? $signed(-32'she610) : $signed(_GEN_694); // @[FFT.scala 35:12]
  assign _GEN_696 = 9'hb7 == cnt[8:0] ? $signed(-32'she6bf) : $signed(_GEN_695); // @[FFT.scala 35:12]
  assign _GEN_697 = 9'hb8 == cnt[8:0] ? $signed(-32'she76c) : $signed(_GEN_696); // @[FFT.scala 35:12]
  assign _GEN_698 = 9'hb9 == cnt[8:0] ? $signed(-32'she817) : $signed(_GEN_697); // @[FFT.scala 35:12]
  assign _GEN_699 = 9'hba == cnt[8:0] ? $signed(-32'she8bf) : $signed(_GEN_698); // @[FFT.scala 35:12]
  assign _GEN_700 = 9'hbb == cnt[8:0] ? $signed(-32'she966) : $signed(_GEN_699); // @[FFT.scala 35:12]
  assign _GEN_701 = 9'hbc == cnt[8:0] ? $signed(-32'shea0a) : $signed(_GEN_700); // @[FFT.scala 35:12]
  assign _GEN_702 = 9'hbd == cnt[8:0] ? $signed(-32'sheaab) : $signed(_GEN_701); // @[FFT.scala 35:12]
  assign _GEN_703 = 9'hbe == cnt[8:0] ? $signed(-32'sheb4b) : $signed(_GEN_702); // @[FFT.scala 35:12]
  assign _GEN_704 = 9'hbf == cnt[8:0] ? $signed(-32'shebe8) : $signed(_GEN_703); // @[FFT.scala 35:12]
  assign _GEN_705 = 9'hc0 == cnt[8:0] ? $signed(-32'shec83) : $signed(_GEN_704); // @[FFT.scala 35:12]
  assign _GEN_706 = 9'hc1 == cnt[8:0] ? $signed(-32'shed1c) : $signed(_GEN_705); // @[FFT.scala 35:12]
  assign _GEN_707 = 9'hc2 == cnt[8:0] ? $signed(-32'shedb3) : $signed(_GEN_706); // @[FFT.scala 35:12]
  assign _GEN_708 = 9'hc3 == cnt[8:0] ? $signed(-32'shee47) : $signed(_GEN_707); // @[FFT.scala 35:12]
  assign _GEN_709 = 9'hc4 == cnt[8:0] ? $signed(-32'sheed9) : $signed(_GEN_708); // @[FFT.scala 35:12]
  assign _GEN_710 = 9'hc5 == cnt[8:0] ? $signed(-32'shef68) : $signed(_GEN_709); // @[FFT.scala 35:12]
  assign _GEN_711 = 9'hc6 == cnt[8:0] ? $signed(-32'sheff5) : $signed(_GEN_710); // @[FFT.scala 35:12]
  assign _GEN_712 = 9'hc7 == cnt[8:0] ? $signed(-32'shf080) : $signed(_GEN_711); // @[FFT.scala 35:12]
  assign _GEN_713 = 9'hc8 == cnt[8:0] ? $signed(-32'shf109) : $signed(_GEN_712); // @[FFT.scala 35:12]
  assign _GEN_714 = 9'hc9 == cnt[8:0] ? $signed(-32'shf18f) : $signed(_GEN_713); // @[FFT.scala 35:12]
  assign _GEN_715 = 9'hca == cnt[8:0] ? $signed(-32'shf213) : $signed(_GEN_714); // @[FFT.scala 35:12]
  assign _GEN_716 = 9'hcb == cnt[8:0] ? $signed(-32'shf295) : $signed(_GEN_715); // @[FFT.scala 35:12]
  assign _GEN_717 = 9'hcc == cnt[8:0] ? $signed(-32'shf314) : $signed(_GEN_716); // @[FFT.scala 35:12]
  assign _GEN_718 = 9'hcd == cnt[8:0] ? $signed(-32'shf391) : $signed(_GEN_717); // @[FFT.scala 35:12]
  assign _GEN_719 = 9'hce == cnt[8:0] ? $signed(-32'shf40c) : $signed(_GEN_718); // @[FFT.scala 35:12]
  assign _GEN_720 = 9'hcf == cnt[8:0] ? $signed(-32'shf484) : $signed(_GEN_719); // @[FFT.scala 35:12]
  assign _GEN_721 = 9'hd0 == cnt[8:0] ? $signed(-32'shf4fa) : $signed(_GEN_720); // @[FFT.scala 35:12]
  assign _GEN_722 = 9'hd1 == cnt[8:0] ? $signed(-32'shf56e) : $signed(_GEN_721); // @[FFT.scala 35:12]
  assign _GEN_723 = 9'hd2 == cnt[8:0] ? $signed(-32'shf5df) : $signed(_GEN_722); // @[FFT.scala 35:12]
  assign _GEN_724 = 9'hd3 == cnt[8:0] ? $signed(-32'shf64e) : $signed(_GEN_723); // @[FFT.scala 35:12]
  assign _GEN_725 = 9'hd4 == cnt[8:0] ? $signed(-32'shf6ba) : $signed(_GEN_724); // @[FFT.scala 35:12]
  assign _GEN_726 = 9'hd5 == cnt[8:0] ? $signed(-32'shf724) : $signed(_GEN_725); // @[FFT.scala 35:12]
  assign _GEN_727 = 9'hd6 == cnt[8:0] ? $signed(-32'shf78c) : $signed(_GEN_726); // @[FFT.scala 35:12]
  assign _GEN_728 = 9'hd7 == cnt[8:0] ? $signed(-32'shf7f1) : $signed(_GEN_727); // @[FFT.scala 35:12]
  assign _GEN_729 = 9'hd8 == cnt[8:0] ? $signed(-32'shf854) : $signed(_GEN_728); // @[FFT.scala 35:12]
  assign _GEN_730 = 9'hd9 == cnt[8:0] ? $signed(-32'shf8b4) : $signed(_GEN_729); // @[FFT.scala 35:12]
  assign _GEN_731 = 9'hda == cnt[8:0] ? $signed(-32'shf913) : $signed(_GEN_730); // @[FFT.scala 35:12]
  assign _GEN_732 = 9'hdb == cnt[8:0] ? $signed(-32'shf96e) : $signed(_GEN_731); // @[FFT.scala 35:12]
  assign _GEN_733 = 9'hdc == cnt[8:0] ? $signed(-32'shf9c8) : $signed(_GEN_732); // @[FFT.scala 35:12]
  assign _GEN_734 = 9'hdd == cnt[8:0] ? $signed(-32'shfa1f) : $signed(_GEN_733); // @[FFT.scala 35:12]
  assign _GEN_735 = 9'hde == cnt[8:0] ? $signed(-32'shfa73) : $signed(_GEN_734); // @[FFT.scala 35:12]
  assign _GEN_736 = 9'hdf == cnt[8:0] ? $signed(-32'shfac5) : $signed(_GEN_735); // @[FFT.scala 35:12]
  assign _GEN_737 = 9'he0 == cnt[8:0] ? $signed(-32'shfb15) : $signed(_GEN_736); // @[FFT.scala 35:12]
  assign _GEN_738 = 9'he1 == cnt[8:0] ? $signed(-32'shfb62) : $signed(_GEN_737); // @[FFT.scala 35:12]
  assign _GEN_739 = 9'he2 == cnt[8:0] ? $signed(-32'shfbad) : $signed(_GEN_738); // @[FFT.scala 35:12]
  assign _GEN_740 = 9'he3 == cnt[8:0] ? $signed(-32'shfbf5) : $signed(_GEN_739); // @[FFT.scala 35:12]
  assign _GEN_741 = 9'he4 == cnt[8:0] ? $signed(-32'shfc3b) : $signed(_GEN_740); // @[FFT.scala 35:12]
  assign _GEN_742 = 9'he5 == cnt[8:0] ? $signed(-32'shfc7f) : $signed(_GEN_741); // @[FFT.scala 35:12]
  assign _GEN_743 = 9'he6 == cnt[8:0] ? $signed(-32'shfcc0) : $signed(_GEN_742); // @[FFT.scala 35:12]
  assign _GEN_744 = 9'he7 == cnt[8:0] ? $signed(-32'shfcfe) : $signed(_GEN_743); // @[FFT.scala 35:12]
  assign _GEN_745 = 9'he8 == cnt[8:0] ? $signed(-32'shfd3b) : $signed(_GEN_744); // @[FFT.scala 35:12]
  assign _GEN_746 = 9'he9 == cnt[8:0] ? $signed(-32'shfd74) : $signed(_GEN_745); // @[FFT.scala 35:12]
  assign _GEN_747 = 9'hea == cnt[8:0] ? $signed(-32'shfdac) : $signed(_GEN_746); // @[FFT.scala 35:12]
  assign _GEN_748 = 9'heb == cnt[8:0] ? $signed(-32'shfde1) : $signed(_GEN_747); // @[FFT.scala 35:12]
  assign _GEN_749 = 9'hec == cnt[8:0] ? $signed(-32'shfe13) : $signed(_GEN_748); // @[FFT.scala 35:12]
  assign _GEN_750 = 9'hed == cnt[8:0] ? $signed(-32'shfe43) : $signed(_GEN_749); // @[FFT.scala 35:12]
  assign _GEN_751 = 9'hee == cnt[8:0] ? $signed(-32'shfe71) : $signed(_GEN_750); // @[FFT.scala 35:12]
  assign _GEN_752 = 9'hef == cnt[8:0] ? $signed(-32'shfe9c) : $signed(_GEN_751); // @[FFT.scala 35:12]
  assign _GEN_753 = 9'hf0 == cnt[8:0] ? $signed(-32'shfec4) : $signed(_GEN_752); // @[FFT.scala 35:12]
  assign _GEN_754 = 9'hf1 == cnt[8:0] ? $signed(-32'shfeeb) : $signed(_GEN_753); // @[FFT.scala 35:12]
  assign _GEN_755 = 9'hf2 == cnt[8:0] ? $signed(-32'shff0e) : $signed(_GEN_754); // @[FFT.scala 35:12]
  assign _GEN_756 = 9'hf3 == cnt[8:0] ? $signed(-32'shff30) : $signed(_GEN_755); // @[FFT.scala 35:12]
  assign _GEN_757 = 9'hf4 == cnt[8:0] ? $signed(-32'shff4e) : $signed(_GEN_756); // @[FFT.scala 35:12]
  assign _GEN_758 = 9'hf5 == cnt[8:0] ? $signed(-32'shff6b) : $signed(_GEN_757); // @[FFT.scala 35:12]
  assign _GEN_759 = 9'hf6 == cnt[8:0] ? $signed(-32'shff85) : $signed(_GEN_758); // @[FFT.scala 35:12]
  assign _GEN_760 = 9'hf7 == cnt[8:0] ? $signed(-32'shff9c) : $signed(_GEN_759); // @[FFT.scala 35:12]
  assign _GEN_761 = 9'hf8 == cnt[8:0] ? $signed(-32'shffb1) : $signed(_GEN_760); // @[FFT.scala 35:12]
  assign _GEN_762 = 9'hf9 == cnt[8:0] ? $signed(-32'shffc4) : $signed(_GEN_761); // @[FFT.scala 35:12]
  assign _GEN_763 = 9'hfa == cnt[8:0] ? $signed(-32'shffd4) : $signed(_GEN_762); // @[FFT.scala 35:12]
  assign _GEN_764 = 9'hfb == cnt[8:0] ? $signed(-32'shffe1) : $signed(_GEN_763); // @[FFT.scala 35:12]
  assign _GEN_765 = 9'hfc == cnt[8:0] ? $signed(-32'shffec) : $signed(_GEN_764); // @[FFT.scala 35:12]
  assign _GEN_766 = 9'hfd == cnt[8:0] ? $signed(-32'shfff5) : $signed(_GEN_765); // @[FFT.scala 35:12]
  assign _GEN_767 = 9'hfe == cnt[8:0] ? $signed(-32'shfffb) : $signed(_GEN_766); // @[FFT.scala 35:12]
  assign _GEN_768 = 9'hff == cnt[8:0] ? $signed(-32'shffff) : $signed(_GEN_767); // @[FFT.scala 35:12]
  assign _GEN_769 = 9'h100 == cnt[8:0] ? $signed(-32'sh10000) : $signed(_GEN_768); // @[FFT.scala 35:12]
  assign _GEN_770 = 9'h101 == cnt[8:0] ? $signed(-32'shffff) : $signed(_GEN_769); // @[FFT.scala 35:12]
  assign _GEN_771 = 9'h102 == cnt[8:0] ? $signed(-32'shfffb) : $signed(_GEN_770); // @[FFT.scala 35:12]
  assign _GEN_772 = 9'h103 == cnt[8:0] ? $signed(-32'shfff5) : $signed(_GEN_771); // @[FFT.scala 35:12]
  assign _GEN_773 = 9'h104 == cnt[8:0] ? $signed(-32'shffec) : $signed(_GEN_772); // @[FFT.scala 35:12]
  assign _GEN_774 = 9'h105 == cnt[8:0] ? $signed(-32'shffe1) : $signed(_GEN_773); // @[FFT.scala 35:12]
  assign _GEN_775 = 9'h106 == cnt[8:0] ? $signed(-32'shffd4) : $signed(_GEN_774); // @[FFT.scala 35:12]
  assign _GEN_776 = 9'h107 == cnt[8:0] ? $signed(-32'shffc4) : $signed(_GEN_775); // @[FFT.scala 35:12]
  assign _GEN_777 = 9'h108 == cnt[8:0] ? $signed(-32'shffb1) : $signed(_GEN_776); // @[FFT.scala 35:12]
  assign _GEN_778 = 9'h109 == cnt[8:0] ? $signed(-32'shff9c) : $signed(_GEN_777); // @[FFT.scala 35:12]
  assign _GEN_779 = 9'h10a == cnt[8:0] ? $signed(-32'shff85) : $signed(_GEN_778); // @[FFT.scala 35:12]
  assign _GEN_780 = 9'h10b == cnt[8:0] ? $signed(-32'shff6b) : $signed(_GEN_779); // @[FFT.scala 35:12]
  assign _GEN_781 = 9'h10c == cnt[8:0] ? $signed(-32'shff4e) : $signed(_GEN_780); // @[FFT.scala 35:12]
  assign _GEN_782 = 9'h10d == cnt[8:0] ? $signed(-32'shff30) : $signed(_GEN_781); // @[FFT.scala 35:12]
  assign _GEN_783 = 9'h10e == cnt[8:0] ? $signed(-32'shff0e) : $signed(_GEN_782); // @[FFT.scala 35:12]
  assign _GEN_784 = 9'h10f == cnt[8:0] ? $signed(-32'shfeeb) : $signed(_GEN_783); // @[FFT.scala 35:12]
  assign _GEN_785 = 9'h110 == cnt[8:0] ? $signed(-32'shfec4) : $signed(_GEN_784); // @[FFT.scala 35:12]
  assign _GEN_786 = 9'h111 == cnt[8:0] ? $signed(-32'shfe9c) : $signed(_GEN_785); // @[FFT.scala 35:12]
  assign _GEN_787 = 9'h112 == cnt[8:0] ? $signed(-32'shfe71) : $signed(_GEN_786); // @[FFT.scala 35:12]
  assign _GEN_788 = 9'h113 == cnt[8:0] ? $signed(-32'shfe43) : $signed(_GEN_787); // @[FFT.scala 35:12]
  assign _GEN_789 = 9'h114 == cnt[8:0] ? $signed(-32'shfe13) : $signed(_GEN_788); // @[FFT.scala 35:12]
  assign _GEN_790 = 9'h115 == cnt[8:0] ? $signed(-32'shfde1) : $signed(_GEN_789); // @[FFT.scala 35:12]
  assign _GEN_791 = 9'h116 == cnt[8:0] ? $signed(-32'shfdac) : $signed(_GEN_790); // @[FFT.scala 35:12]
  assign _GEN_792 = 9'h117 == cnt[8:0] ? $signed(-32'shfd74) : $signed(_GEN_791); // @[FFT.scala 35:12]
  assign _GEN_793 = 9'h118 == cnt[8:0] ? $signed(-32'shfd3b) : $signed(_GEN_792); // @[FFT.scala 35:12]
  assign _GEN_794 = 9'h119 == cnt[8:0] ? $signed(-32'shfcfe) : $signed(_GEN_793); // @[FFT.scala 35:12]
  assign _GEN_795 = 9'h11a == cnt[8:0] ? $signed(-32'shfcc0) : $signed(_GEN_794); // @[FFT.scala 35:12]
  assign _GEN_796 = 9'h11b == cnt[8:0] ? $signed(-32'shfc7f) : $signed(_GEN_795); // @[FFT.scala 35:12]
  assign _GEN_797 = 9'h11c == cnt[8:0] ? $signed(-32'shfc3b) : $signed(_GEN_796); // @[FFT.scala 35:12]
  assign _GEN_798 = 9'h11d == cnt[8:0] ? $signed(-32'shfbf5) : $signed(_GEN_797); // @[FFT.scala 35:12]
  assign _GEN_799 = 9'h11e == cnt[8:0] ? $signed(-32'shfbad) : $signed(_GEN_798); // @[FFT.scala 35:12]
  assign _GEN_800 = 9'h11f == cnt[8:0] ? $signed(-32'shfb62) : $signed(_GEN_799); // @[FFT.scala 35:12]
  assign _GEN_801 = 9'h120 == cnt[8:0] ? $signed(-32'shfb15) : $signed(_GEN_800); // @[FFT.scala 35:12]
  assign _GEN_802 = 9'h121 == cnt[8:0] ? $signed(-32'shfac5) : $signed(_GEN_801); // @[FFT.scala 35:12]
  assign _GEN_803 = 9'h122 == cnt[8:0] ? $signed(-32'shfa73) : $signed(_GEN_802); // @[FFT.scala 35:12]
  assign _GEN_804 = 9'h123 == cnt[8:0] ? $signed(-32'shfa1f) : $signed(_GEN_803); // @[FFT.scala 35:12]
  assign _GEN_805 = 9'h124 == cnt[8:0] ? $signed(-32'shf9c8) : $signed(_GEN_804); // @[FFT.scala 35:12]
  assign _GEN_806 = 9'h125 == cnt[8:0] ? $signed(-32'shf96e) : $signed(_GEN_805); // @[FFT.scala 35:12]
  assign _GEN_807 = 9'h126 == cnt[8:0] ? $signed(-32'shf913) : $signed(_GEN_806); // @[FFT.scala 35:12]
  assign _GEN_808 = 9'h127 == cnt[8:0] ? $signed(-32'shf8b4) : $signed(_GEN_807); // @[FFT.scala 35:12]
  assign _GEN_809 = 9'h128 == cnt[8:0] ? $signed(-32'shf854) : $signed(_GEN_808); // @[FFT.scala 35:12]
  assign _GEN_810 = 9'h129 == cnt[8:0] ? $signed(-32'shf7f1) : $signed(_GEN_809); // @[FFT.scala 35:12]
  assign _GEN_811 = 9'h12a == cnt[8:0] ? $signed(-32'shf78c) : $signed(_GEN_810); // @[FFT.scala 35:12]
  assign _GEN_812 = 9'h12b == cnt[8:0] ? $signed(-32'shf724) : $signed(_GEN_811); // @[FFT.scala 35:12]
  assign _GEN_813 = 9'h12c == cnt[8:0] ? $signed(-32'shf6ba) : $signed(_GEN_812); // @[FFT.scala 35:12]
  assign _GEN_814 = 9'h12d == cnt[8:0] ? $signed(-32'shf64e) : $signed(_GEN_813); // @[FFT.scala 35:12]
  assign _GEN_815 = 9'h12e == cnt[8:0] ? $signed(-32'shf5df) : $signed(_GEN_814); // @[FFT.scala 35:12]
  assign _GEN_816 = 9'h12f == cnt[8:0] ? $signed(-32'shf56e) : $signed(_GEN_815); // @[FFT.scala 35:12]
  assign _GEN_817 = 9'h130 == cnt[8:0] ? $signed(-32'shf4fa) : $signed(_GEN_816); // @[FFT.scala 35:12]
  assign _GEN_818 = 9'h131 == cnt[8:0] ? $signed(-32'shf484) : $signed(_GEN_817); // @[FFT.scala 35:12]
  assign _GEN_819 = 9'h132 == cnt[8:0] ? $signed(-32'shf40c) : $signed(_GEN_818); // @[FFT.scala 35:12]
  assign _GEN_820 = 9'h133 == cnt[8:0] ? $signed(-32'shf391) : $signed(_GEN_819); // @[FFT.scala 35:12]
  assign _GEN_821 = 9'h134 == cnt[8:0] ? $signed(-32'shf314) : $signed(_GEN_820); // @[FFT.scala 35:12]
  assign _GEN_822 = 9'h135 == cnt[8:0] ? $signed(-32'shf295) : $signed(_GEN_821); // @[FFT.scala 35:12]
  assign _GEN_823 = 9'h136 == cnt[8:0] ? $signed(-32'shf213) : $signed(_GEN_822); // @[FFT.scala 35:12]
  assign _GEN_824 = 9'h137 == cnt[8:0] ? $signed(-32'shf18f) : $signed(_GEN_823); // @[FFT.scala 35:12]
  assign _GEN_825 = 9'h138 == cnt[8:0] ? $signed(-32'shf109) : $signed(_GEN_824); // @[FFT.scala 35:12]
  assign _GEN_826 = 9'h139 == cnt[8:0] ? $signed(-32'shf080) : $signed(_GEN_825); // @[FFT.scala 35:12]
  assign _GEN_827 = 9'h13a == cnt[8:0] ? $signed(-32'sheff5) : $signed(_GEN_826); // @[FFT.scala 35:12]
  assign _GEN_828 = 9'h13b == cnt[8:0] ? $signed(-32'shef68) : $signed(_GEN_827); // @[FFT.scala 35:12]
  assign _GEN_829 = 9'h13c == cnt[8:0] ? $signed(-32'sheed9) : $signed(_GEN_828); // @[FFT.scala 35:12]
  assign _GEN_830 = 9'h13d == cnt[8:0] ? $signed(-32'shee47) : $signed(_GEN_829); // @[FFT.scala 35:12]
  assign _GEN_831 = 9'h13e == cnt[8:0] ? $signed(-32'shedb3) : $signed(_GEN_830); // @[FFT.scala 35:12]
  assign _GEN_832 = 9'h13f == cnt[8:0] ? $signed(-32'shed1c) : $signed(_GEN_831); // @[FFT.scala 35:12]
  assign _GEN_833 = 9'h140 == cnt[8:0] ? $signed(-32'shec83) : $signed(_GEN_832); // @[FFT.scala 35:12]
  assign _GEN_834 = 9'h141 == cnt[8:0] ? $signed(-32'shebe8) : $signed(_GEN_833); // @[FFT.scala 35:12]
  assign _GEN_835 = 9'h142 == cnt[8:0] ? $signed(-32'sheb4b) : $signed(_GEN_834); // @[FFT.scala 35:12]
  assign _GEN_836 = 9'h143 == cnt[8:0] ? $signed(-32'sheaab) : $signed(_GEN_835); // @[FFT.scala 35:12]
  assign _GEN_837 = 9'h144 == cnt[8:0] ? $signed(-32'shea0a) : $signed(_GEN_836); // @[FFT.scala 35:12]
  assign _GEN_838 = 9'h145 == cnt[8:0] ? $signed(-32'she966) : $signed(_GEN_837); // @[FFT.scala 35:12]
  assign _GEN_839 = 9'h146 == cnt[8:0] ? $signed(-32'she8bf) : $signed(_GEN_838); // @[FFT.scala 35:12]
  assign _GEN_840 = 9'h147 == cnt[8:0] ? $signed(-32'she817) : $signed(_GEN_839); // @[FFT.scala 35:12]
  assign _GEN_841 = 9'h148 == cnt[8:0] ? $signed(-32'she76c) : $signed(_GEN_840); // @[FFT.scala 35:12]
  assign _GEN_842 = 9'h149 == cnt[8:0] ? $signed(-32'she6bf) : $signed(_GEN_841); // @[FFT.scala 35:12]
  assign _GEN_843 = 9'h14a == cnt[8:0] ? $signed(-32'she610) : $signed(_GEN_842); // @[FFT.scala 35:12]
  assign _GEN_844 = 9'h14b == cnt[8:0] ? $signed(-32'she55e) : $signed(_GEN_843); // @[FFT.scala 35:12]
  assign _GEN_845 = 9'h14c == cnt[8:0] ? $signed(-32'she4aa) : $signed(_GEN_844); // @[FFT.scala 35:12]
  assign _GEN_846 = 9'h14d == cnt[8:0] ? $signed(-32'she3f4) : $signed(_GEN_845); // @[FFT.scala 35:12]
  assign _GEN_847 = 9'h14e == cnt[8:0] ? $signed(-32'she33c) : $signed(_GEN_846); // @[FFT.scala 35:12]
  assign _GEN_848 = 9'h14f == cnt[8:0] ? $signed(-32'she282) : $signed(_GEN_847); // @[FFT.scala 35:12]
  assign _GEN_849 = 9'h150 == cnt[8:0] ? $signed(-32'she1c6) : $signed(_GEN_848); // @[FFT.scala 35:12]
  assign _GEN_850 = 9'h151 == cnt[8:0] ? $signed(-32'she107) : $signed(_GEN_849); // @[FFT.scala 35:12]
  assign _GEN_851 = 9'h152 == cnt[8:0] ? $signed(-32'she046) : $signed(_GEN_850); // @[FFT.scala 35:12]
  assign _GEN_852 = 9'h153 == cnt[8:0] ? $signed(-32'shdf83) : $signed(_GEN_851); // @[FFT.scala 35:12]
  assign _GEN_853 = 9'h154 == cnt[8:0] ? $signed(-32'shdebe) : $signed(_GEN_852); // @[FFT.scala 35:12]
  assign _GEN_854 = 9'h155 == cnt[8:0] ? $signed(-32'shddf7) : $signed(_GEN_853); // @[FFT.scala 35:12]
  assign _GEN_855 = 9'h156 == cnt[8:0] ? $signed(-32'shdd2d) : $signed(_GEN_854); // @[FFT.scala 35:12]
  assign _GEN_856 = 9'h157 == cnt[8:0] ? $signed(-32'shdc62) : $signed(_GEN_855); // @[FFT.scala 35:12]
  assign _GEN_857 = 9'h158 == cnt[8:0] ? $signed(-32'shdb94) : $signed(_GEN_856); // @[FFT.scala 35:12]
  assign _GEN_858 = 9'h159 == cnt[8:0] ? $signed(-32'shdac4) : $signed(_GEN_857); // @[FFT.scala 35:12]
  assign _GEN_859 = 9'h15a == cnt[8:0] ? $signed(-32'shd9f2) : $signed(_GEN_858); // @[FFT.scala 35:12]
  assign _GEN_860 = 9'h15b == cnt[8:0] ? $signed(-32'shd91e) : $signed(_GEN_859); // @[FFT.scala 35:12]
  assign _GEN_861 = 9'h15c == cnt[8:0] ? $signed(-32'shd848) : $signed(_GEN_860); // @[FFT.scala 35:12]
  assign _GEN_862 = 9'h15d == cnt[8:0] ? $signed(-32'shd770) : $signed(_GEN_861); // @[FFT.scala 35:12]
  assign _GEN_863 = 9'h15e == cnt[8:0] ? $signed(-32'shd696) : $signed(_GEN_862); // @[FFT.scala 35:12]
  assign _GEN_864 = 9'h15f == cnt[8:0] ? $signed(-32'shd5ba) : $signed(_GEN_863); // @[FFT.scala 35:12]
  assign _GEN_865 = 9'h160 == cnt[8:0] ? $signed(-32'shd4db) : $signed(_GEN_864); // @[FFT.scala 35:12]
  assign _GEN_866 = 9'h161 == cnt[8:0] ? $signed(-32'shd3fb) : $signed(_GEN_865); // @[FFT.scala 35:12]
  assign _GEN_867 = 9'h162 == cnt[8:0] ? $signed(-32'shd318) : $signed(_GEN_866); // @[FFT.scala 35:12]
  assign _GEN_868 = 9'h163 == cnt[8:0] ? $signed(-32'shd234) : $signed(_GEN_867); // @[FFT.scala 35:12]
  assign _GEN_869 = 9'h164 == cnt[8:0] ? $signed(-32'shd14d) : $signed(_GEN_868); // @[FFT.scala 35:12]
  assign _GEN_870 = 9'h165 == cnt[8:0] ? $signed(-32'shd065) : $signed(_GEN_869); // @[FFT.scala 35:12]
  assign _GEN_871 = 9'h166 == cnt[8:0] ? $signed(-32'shcf7a) : $signed(_GEN_870); // @[FFT.scala 35:12]
  assign _GEN_872 = 9'h167 == cnt[8:0] ? $signed(-32'shce8e) : $signed(_GEN_871); // @[FFT.scala 35:12]
  assign _GEN_873 = 9'h168 == cnt[8:0] ? $signed(-32'shcd9f) : $signed(_GEN_872); // @[FFT.scala 35:12]
  assign _GEN_874 = 9'h169 == cnt[8:0] ? $signed(-32'shccae) : $signed(_GEN_873); // @[FFT.scala 35:12]
  assign _GEN_875 = 9'h16a == cnt[8:0] ? $signed(-32'shcbbc) : $signed(_GEN_874); // @[FFT.scala 35:12]
  assign _GEN_876 = 9'h16b == cnt[8:0] ? $signed(-32'shcac7) : $signed(_GEN_875); // @[FFT.scala 35:12]
  assign _GEN_877 = 9'h16c == cnt[8:0] ? $signed(-32'shc9d1) : $signed(_GEN_876); // @[FFT.scala 35:12]
  assign _GEN_878 = 9'h16d == cnt[8:0] ? $signed(-32'shc8d9) : $signed(_GEN_877); // @[FFT.scala 35:12]
  assign _GEN_879 = 9'h16e == cnt[8:0] ? $signed(-32'shc7de) : $signed(_GEN_878); // @[FFT.scala 35:12]
  assign _GEN_880 = 9'h16f == cnt[8:0] ? $signed(-32'shc6e2) : $signed(_GEN_879); // @[FFT.scala 35:12]
  assign _GEN_881 = 9'h170 == cnt[8:0] ? $signed(-32'shc5e4) : $signed(_GEN_880); // @[FFT.scala 35:12]
  assign _GEN_882 = 9'h171 == cnt[8:0] ? $signed(-32'shc4e4) : $signed(_GEN_881); // @[FFT.scala 35:12]
  assign _GEN_883 = 9'h172 == cnt[8:0] ? $signed(-32'shc3e2) : $signed(_GEN_882); // @[FFT.scala 35:12]
  assign _GEN_884 = 9'h173 == cnt[8:0] ? $signed(-32'shc2de) : $signed(_GEN_883); // @[FFT.scala 35:12]
  assign _GEN_885 = 9'h174 == cnt[8:0] ? $signed(-32'shc1d8) : $signed(_GEN_884); // @[FFT.scala 35:12]
  assign _GEN_886 = 9'h175 == cnt[8:0] ? $signed(-32'shc0d1) : $signed(_GEN_885); // @[FFT.scala 35:12]
  assign _GEN_887 = 9'h176 == cnt[8:0] ? $signed(-32'shbfc7) : $signed(_GEN_886); // @[FFT.scala 35:12]
  assign _GEN_888 = 9'h177 == cnt[8:0] ? $signed(-32'shbebc) : $signed(_GEN_887); // @[FFT.scala 35:12]
  assign _GEN_889 = 9'h178 == cnt[8:0] ? $signed(-32'shbdaf) : $signed(_GEN_888); // @[FFT.scala 35:12]
  assign _GEN_890 = 9'h179 == cnt[8:0] ? $signed(-32'shbca0) : $signed(_GEN_889); // @[FFT.scala 35:12]
  assign _GEN_891 = 9'h17a == cnt[8:0] ? $signed(-32'shbb8f) : $signed(_GEN_890); // @[FFT.scala 35:12]
  assign _GEN_892 = 9'h17b == cnt[8:0] ? $signed(-32'shba7d) : $signed(_GEN_891); // @[FFT.scala 35:12]
  assign _GEN_893 = 9'h17c == cnt[8:0] ? $signed(-32'shb968) : $signed(_GEN_892); // @[FFT.scala 35:12]
  assign _GEN_894 = 9'h17d == cnt[8:0] ? $signed(-32'shb852) : $signed(_GEN_893); // @[FFT.scala 35:12]
  assign _GEN_895 = 9'h17e == cnt[8:0] ? $signed(-32'shb73a) : $signed(_GEN_894); // @[FFT.scala 35:12]
  assign _GEN_896 = 9'h17f == cnt[8:0] ? $signed(-32'shb620) : $signed(_GEN_895); // @[FFT.scala 35:12]
  assign _GEN_897 = 9'h180 == cnt[8:0] ? $signed(-32'shb505) : $signed(_GEN_896); // @[FFT.scala 35:12]
  assign _GEN_898 = 9'h181 == cnt[8:0] ? $signed(-32'shb3e8) : $signed(_GEN_897); // @[FFT.scala 35:12]
  assign _GEN_899 = 9'h182 == cnt[8:0] ? $signed(-32'shb2c9) : $signed(_GEN_898); // @[FFT.scala 35:12]
  assign _GEN_900 = 9'h183 == cnt[8:0] ? $signed(-32'shb1a8) : $signed(_GEN_899); // @[FFT.scala 35:12]
  assign _GEN_901 = 9'h184 == cnt[8:0] ? $signed(-32'shb086) : $signed(_GEN_900); // @[FFT.scala 35:12]
  assign _GEN_902 = 9'h185 == cnt[8:0] ? $signed(-32'shaf62) : $signed(_GEN_901); // @[FFT.scala 35:12]
  assign _GEN_903 = 9'h186 == cnt[8:0] ? $signed(-32'shae3c) : $signed(_GEN_902); // @[FFT.scala 35:12]
  assign _GEN_904 = 9'h187 == cnt[8:0] ? $signed(-32'shad14) : $signed(_GEN_903); // @[FFT.scala 35:12]
  assign _GEN_905 = 9'h188 == cnt[8:0] ? $signed(-32'shabeb) : $signed(_GEN_904); // @[FFT.scala 35:12]
  assign _GEN_906 = 9'h189 == cnt[8:0] ? $signed(-32'shaac1) : $signed(_GEN_905); // @[FFT.scala 35:12]
  assign _GEN_907 = 9'h18a == cnt[8:0] ? $signed(-32'sha994) : $signed(_GEN_906); // @[FFT.scala 35:12]
  assign _GEN_908 = 9'h18b == cnt[8:0] ? $signed(-32'sha866) : $signed(_GEN_907); // @[FFT.scala 35:12]
  assign _GEN_909 = 9'h18c == cnt[8:0] ? $signed(-32'sha736) : $signed(_GEN_908); // @[FFT.scala 35:12]
  assign _GEN_910 = 9'h18d == cnt[8:0] ? $signed(-32'sha605) : $signed(_GEN_909); // @[FFT.scala 35:12]
  assign _GEN_911 = 9'h18e == cnt[8:0] ? $signed(-32'sha4d2) : $signed(_GEN_910); // @[FFT.scala 35:12]
  assign _GEN_912 = 9'h18f == cnt[8:0] ? $signed(-32'sha39e) : $signed(_GEN_911); // @[FFT.scala 35:12]
  assign _GEN_913 = 9'h190 == cnt[8:0] ? $signed(-32'sha268) : $signed(_GEN_912); // @[FFT.scala 35:12]
  assign _GEN_914 = 9'h191 == cnt[8:0] ? $signed(-32'sha130) : $signed(_GEN_913); // @[FFT.scala 35:12]
  assign _GEN_915 = 9'h192 == cnt[8:0] ? $signed(-32'sh9ff7) : $signed(_GEN_914); // @[FFT.scala 35:12]
  assign _GEN_916 = 9'h193 == cnt[8:0] ? $signed(-32'sh9ebc) : $signed(_GEN_915); // @[FFT.scala 35:12]
  assign _GEN_917 = 9'h194 == cnt[8:0] ? $signed(-32'sh9d80) : $signed(_GEN_916); // @[FFT.scala 35:12]
  assign _GEN_918 = 9'h195 == cnt[8:0] ? $signed(-32'sh9c42) : $signed(_GEN_917); // @[FFT.scala 35:12]
  assign _GEN_919 = 9'h196 == cnt[8:0] ? $signed(-32'sh9b03) : $signed(_GEN_918); // @[FFT.scala 35:12]
  assign _GEN_920 = 9'h197 == cnt[8:0] ? $signed(-32'sh99c2) : $signed(_GEN_919); // @[FFT.scala 35:12]
  assign _GEN_921 = 9'h198 == cnt[8:0] ? $signed(-32'sh9880) : $signed(_GEN_920); // @[FFT.scala 35:12]
  assign _GEN_922 = 9'h199 == cnt[8:0] ? $signed(-32'sh973c) : $signed(_GEN_921); // @[FFT.scala 35:12]
  assign _GEN_923 = 9'h19a == cnt[8:0] ? $signed(-32'sh95f7) : $signed(_GEN_922); // @[FFT.scala 35:12]
  assign _GEN_924 = 9'h19b == cnt[8:0] ? $signed(-32'sh94b0) : $signed(_GEN_923); // @[FFT.scala 35:12]
  assign _GEN_925 = 9'h19c == cnt[8:0] ? $signed(-32'sh9368) : $signed(_GEN_924); // @[FFT.scala 35:12]
  assign _GEN_926 = 9'h19d == cnt[8:0] ? $signed(-32'sh921f) : $signed(_GEN_925); // @[FFT.scala 35:12]
  assign _GEN_927 = 9'h19e == cnt[8:0] ? $signed(-32'sh90d4) : $signed(_GEN_926); // @[FFT.scala 35:12]
  assign _GEN_928 = 9'h19f == cnt[8:0] ? $signed(-32'sh8f88) : $signed(_GEN_927); // @[FFT.scala 35:12]
  assign _GEN_929 = 9'h1a0 == cnt[8:0] ? $signed(-32'sh8e3a) : $signed(_GEN_928); // @[FFT.scala 35:12]
  assign _GEN_930 = 9'h1a1 == cnt[8:0] ? $signed(-32'sh8ceb) : $signed(_GEN_929); // @[FFT.scala 35:12]
  assign _GEN_931 = 9'h1a2 == cnt[8:0] ? $signed(-32'sh8b9a) : $signed(_GEN_930); // @[FFT.scala 35:12]
  assign _GEN_932 = 9'h1a3 == cnt[8:0] ? $signed(-32'sh8a49) : $signed(_GEN_931); // @[FFT.scala 35:12]
  assign _GEN_933 = 9'h1a4 == cnt[8:0] ? $signed(-32'sh88f6) : $signed(_GEN_932); // @[FFT.scala 35:12]
  assign _GEN_934 = 9'h1a5 == cnt[8:0] ? $signed(-32'sh87a1) : $signed(_GEN_933); // @[FFT.scala 35:12]
  assign _GEN_935 = 9'h1a6 == cnt[8:0] ? $signed(-32'sh864c) : $signed(_GEN_934); // @[FFT.scala 35:12]
  assign _GEN_936 = 9'h1a7 == cnt[8:0] ? $signed(-32'sh84f5) : $signed(_GEN_935); // @[FFT.scala 35:12]
  assign _GEN_937 = 9'h1a8 == cnt[8:0] ? $signed(-32'sh839c) : $signed(_GEN_936); // @[FFT.scala 35:12]
  assign _GEN_938 = 9'h1a9 == cnt[8:0] ? $signed(-32'sh8243) : $signed(_GEN_937); // @[FFT.scala 35:12]
  assign _GEN_939 = 9'h1aa == cnt[8:0] ? $signed(-32'sh80e8) : $signed(_GEN_938); // @[FFT.scala 35:12]
  assign _GEN_940 = 9'h1ab == cnt[8:0] ? $signed(-32'sh7f8c) : $signed(_GEN_939); // @[FFT.scala 35:12]
  assign _GEN_941 = 9'h1ac == cnt[8:0] ? $signed(-32'sh7e2f) : $signed(_GEN_940); // @[FFT.scala 35:12]
  assign _GEN_942 = 9'h1ad == cnt[8:0] ? $signed(-32'sh7cd0) : $signed(_GEN_941); // @[FFT.scala 35:12]
  assign _GEN_943 = 9'h1ae == cnt[8:0] ? $signed(-32'sh7b70) : $signed(_GEN_942); // @[FFT.scala 35:12]
  assign _GEN_944 = 9'h1af == cnt[8:0] ? $signed(-32'sh7a10) : $signed(_GEN_943); // @[FFT.scala 35:12]
  assign _GEN_945 = 9'h1b0 == cnt[8:0] ? $signed(-32'sh78ad) : $signed(_GEN_944); // @[FFT.scala 35:12]
  assign _GEN_946 = 9'h1b1 == cnt[8:0] ? $signed(-32'sh774a) : $signed(_GEN_945); // @[FFT.scala 35:12]
  assign _GEN_947 = 9'h1b2 == cnt[8:0] ? $signed(-32'sh75e6) : $signed(_GEN_946); // @[FFT.scala 35:12]
  assign _GEN_948 = 9'h1b3 == cnt[8:0] ? $signed(-32'sh7480) : $signed(_GEN_947); // @[FFT.scala 35:12]
  assign _GEN_949 = 9'h1b4 == cnt[8:0] ? $signed(-32'sh731a) : $signed(_GEN_948); // @[FFT.scala 35:12]
  assign _GEN_950 = 9'h1b5 == cnt[8:0] ? $signed(-32'sh71b2) : $signed(_GEN_949); // @[FFT.scala 35:12]
  assign _GEN_951 = 9'h1b6 == cnt[8:0] ? $signed(-32'sh7049) : $signed(_GEN_950); // @[FFT.scala 35:12]
  assign _GEN_952 = 9'h1b7 == cnt[8:0] ? $signed(-32'sh6edf) : $signed(_GEN_951); // @[FFT.scala 35:12]
  assign _GEN_953 = 9'h1b8 == cnt[8:0] ? $signed(-32'sh6d74) : $signed(_GEN_952); // @[FFT.scala 35:12]
  assign _GEN_954 = 9'h1b9 == cnt[8:0] ? $signed(-32'sh6c08) : $signed(_GEN_953); // @[FFT.scala 35:12]
  assign _GEN_955 = 9'h1ba == cnt[8:0] ? $signed(-32'sh6a9b) : $signed(_GEN_954); // @[FFT.scala 35:12]
  assign _GEN_956 = 9'h1bb == cnt[8:0] ? $signed(-32'sh692d) : $signed(_GEN_955); // @[FFT.scala 35:12]
  assign _GEN_957 = 9'h1bc == cnt[8:0] ? $signed(-32'sh67be) : $signed(_GEN_956); // @[FFT.scala 35:12]
  assign _GEN_958 = 9'h1bd == cnt[8:0] ? $signed(-32'sh664e) : $signed(_GEN_957); // @[FFT.scala 35:12]
  assign _GEN_959 = 9'h1be == cnt[8:0] ? $signed(-32'sh64dd) : $signed(_GEN_958); // @[FFT.scala 35:12]
  assign _GEN_960 = 9'h1bf == cnt[8:0] ? $signed(-32'sh636b) : $signed(_GEN_959); // @[FFT.scala 35:12]
  assign _GEN_961 = 9'h1c0 == cnt[8:0] ? $signed(-32'sh61f8) : $signed(_GEN_960); // @[FFT.scala 35:12]
  assign _GEN_962 = 9'h1c1 == cnt[8:0] ? $signed(-32'sh6084) : $signed(_GEN_961); // @[FFT.scala 35:12]
  assign _GEN_963 = 9'h1c2 == cnt[8:0] ? $signed(-32'sh5f0f) : $signed(_GEN_962); // @[FFT.scala 35:12]
  assign _GEN_964 = 9'h1c3 == cnt[8:0] ? $signed(-32'sh5d99) : $signed(_GEN_963); // @[FFT.scala 35:12]
  assign _GEN_965 = 9'h1c4 == cnt[8:0] ? $signed(-32'sh5c22) : $signed(_GEN_964); // @[FFT.scala 35:12]
  assign _GEN_966 = 9'h1c5 == cnt[8:0] ? $signed(-32'sh5aaa) : $signed(_GEN_965); // @[FFT.scala 35:12]
  assign _GEN_967 = 9'h1c6 == cnt[8:0] ? $signed(-32'sh5932) : $signed(_GEN_966); // @[FFT.scala 35:12]
  assign _GEN_968 = 9'h1c7 == cnt[8:0] ? $signed(-32'sh57b9) : $signed(_GEN_967); // @[FFT.scala 35:12]
  assign _GEN_969 = 9'h1c8 == cnt[8:0] ? $signed(-32'sh563e) : $signed(_GEN_968); // @[FFT.scala 35:12]
  assign _GEN_970 = 9'h1c9 == cnt[8:0] ? $signed(-32'sh54c3) : $signed(_GEN_969); // @[FFT.scala 35:12]
  assign _GEN_971 = 9'h1ca == cnt[8:0] ? $signed(-32'sh5348) : $signed(_GEN_970); // @[FFT.scala 35:12]
  assign _GEN_972 = 9'h1cb == cnt[8:0] ? $signed(-32'sh51cb) : $signed(_GEN_971); // @[FFT.scala 35:12]
  assign _GEN_973 = 9'h1cc == cnt[8:0] ? $signed(-32'sh504d) : $signed(_GEN_972); // @[FFT.scala 35:12]
  assign _GEN_974 = 9'h1cd == cnt[8:0] ? $signed(-32'sh4ecf) : $signed(_GEN_973); // @[FFT.scala 35:12]
  assign _GEN_975 = 9'h1ce == cnt[8:0] ? $signed(-32'sh4d50) : $signed(_GEN_974); // @[FFT.scala 35:12]
  assign _GEN_976 = 9'h1cf == cnt[8:0] ? $signed(-32'sh4bd1) : $signed(_GEN_975); // @[FFT.scala 35:12]
  assign _GEN_977 = 9'h1d0 == cnt[8:0] ? $signed(-32'sh4a50) : $signed(_GEN_976); // @[FFT.scala 35:12]
  assign _GEN_978 = 9'h1d1 == cnt[8:0] ? $signed(-32'sh48cf) : $signed(_GEN_977); // @[FFT.scala 35:12]
  assign _GEN_979 = 9'h1d2 == cnt[8:0] ? $signed(-32'sh474d) : $signed(_GEN_978); // @[FFT.scala 35:12]
  assign _GEN_980 = 9'h1d3 == cnt[8:0] ? $signed(-32'sh45cb) : $signed(_GEN_979); // @[FFT.scala 35:12]
  assign _GEN_981 = 9'h1d4 == cnt[8:0] ? $signed(-32'sh4447) : $signed(_GEN_980); // @[FFT.scala 35:12]
  assign _GEN_982 = 9'h1d5 == cnt[8:0] ? $signed(-32'sh42c3) : $signed(_GEN_981); // @[FFT.scala 35:12]
  assign _GEN_983 = 9'h1d6 == cnt[8:0] ? $signed(-32'sh413f) : $signed(_GEN_982); // @[FFT.scala 35:12]
  assign _GEN_984 = 9'h1d7 == cnt[8:0] ? $signed(-32'sh3fba) : $signed(_GEN_983); // @[FFT.scala 35:12]
  assign _GEN_985 = 9'h1d8 == cnt[8:0] ? $signed(-32'sh3e34) : $signed(_GEN_984); // @[FFT.scala 35:12]
  assign _GEN_986 = 9'h1d9 == cnt[8:0] ? $signed(-32'sh3cae) : $signed(_GEN_985); // @[FFT.scala 35:12]
  assign _GEN_987 = 9'h1da == cnt[8:0] ? $signed(-32'sh3b27) : $signed(_GEN_986); // @[FFT.scala 35:12]
  assign _GEN_988 = 9'h1db == cnt[8:0] ? $signed(-32'sh399f) : $signed(_GEN_987); // @[FFT.scala 35:12]
  assign _GEN_989 = 9'h1dc == cnt[8:0] ? $signed(-32'sh3817) : $signed(_GEN_988); // @[FFT.scala 35:12]
  assign _GEN_990 = 9'h1dd == cnt[8:0] ? $signed(-32'sh368e) : $signed(_GEN_989); // @[FFT.scala 35:12]
  assign _GEN_991 = 9'h1de == cnt[8:0] ? $signed(-32'sh3505) : $signed(_GEN_990); // @[FFT.scala 35:12]
  assign _GEN_992 = 9'h1df == cnt[8:0] ? $signed(-32'sh337c) : $signed(_GEN_991); // @[FFT.scala 35:12]
  assign _GEN_993 = 9'h1e0 == cnt[8:0] ? $signed(-32'sh31f1) : $signed(_GEN_992); // @[FFT.scala 35:12]
  assign _GEN_994 = 9'h1e1 == cnt[8:0] ? $signed(-32'sh3067) : $signed(_GEN_993); // @[FFT.scala 35:12]
  assign _GEN_995 = 9'h1e2 == cnt[8:0] ? $signed(-32'sh2edc) : $signed(_GEN_994); // @[FFT.scala 35:12]
  assign _GEN_996 = 9'h1e3 == cnt[8:0] ? $signed(-32'sh2d50) : $signed(_GEN_995); // @[FFT.scala 35:12]
  assign _GEN_997 = 9'h1e4 == cnt[8:0] ? $signed(-32'sh2bc4) : $signed(_GEN_996); // @[FFT.scala 35:12]
  assign _GEN_998 = 9'h1e5 == cnt[8:0] ? $signed(-32'sh2a38) : $signed(_GEN_997); // @[FFT.scala 35:12]
  assign _GEN_999 = 9'h1e6 == cnt[8:0] ? $signed(-32'sh28ab) : $signed(_GEN_998); // @[FFT.scala 35:12]
  assign _GEN_1000 = 9'h1e7 == cnt[8:0] ? $signed(-32'sh271e) : $signed(_GEN_999); // @[FFT.scala 35:12]
  assign _GEN_1001 = 9'h1e8 == cnt[8:0] ? $signed(-32'sh2590) : $signed(_GEN_1000); // @[FFT.scala 35:12]
  assign _GEN_1002 = 9'h1e9 == cnt[8:0] ? $signed(-32'sh2402) : $signed(_GEN_1001); // @[FFT.scala 35:12]
  assign _GEN_1003 = 9'h1ea == cnt[8:0] ? $signed(-32'sh2274) : $signed(_GEN_1002); // @[FFT.scala 35:12]
  assign _GEN_1004 = 9'h1eb == cnt[8:0] ? $signed(-32'sh20e5) : $signed(_GEN_1003); // @[FFT.scala 35:12]
  assign _GEN_1005 = 9'h1ec == cnt[8:0] ? $signed(-32'sh1f56) : $signed(_GEN_1004); // @[FFT.scala 35:12]
  assign _GEN_1006 = 9'h1ed == cnt[8:0] ? $signed(-32'sh1dc7) : $signed(_GEN_1005); // @[FFT.scala 35:12]
  assign _GEN_1007 = 9'h1ee == cnt[8:0] ? $signed(-32'sh1c38) : $signed(_GEN_1006); // @[FFT.scala 35:12]
  assign _GEN_1008 = 9'h1ef == cnt[8:0] ? $signed(-32'sh1aa8) : $signed(_GEN_1007); // @[FFT.scala 35:12]
  assign _GEN_1009 = 9'h1f0 == cnt[8:0] ? $signed(-32'sh1918) : $signed(_GEN_1008); // @[FFT.scala 35:12]
  assign _GEN_1010 = 9'h1f1 == cnt[8:0] ? $signed(-32'sh1787) : $signed(_GEN_1009); // @[FFT.scala 35:12]
  assign _GEN_1011 = 9'h1f2 == cnt[8:0] ? $signed(-32'sh15f7) : $signed(_GEN_1010); // @[FFT.scala 35:12]
  assign _GEN_1012 = 9'h1f3 == cnt[8:0] ? $signed(-32'sh1466) : $signed(_GEN_1011); // @[FFT.scala 35:12]
  assign _GEN_1013 = 9'h1f4 == cnt[8:0] ? $signed(-32'sh12d5) : $signed(_GEN_1012); // @[FFT.scala 35:12]
  assign _GEN_1014 = 9'h1f5 == cnt[8:0] ? $signed(-32'sh1144) : $signed(_GEN_1013); // @[FFT.scala 35:12]
  assign _GEN_1015 = 9'h1f6 == cnt[8:0] ? $signed(-32'shfb3) : $signed(_GEN_1014); // @[FFT.scala 35:12]
  assign _GEN_1016 = 9'h1f7 == cnt[8:0] ? $signed(-32'she21) : $signed(_GEN_1015); // @[FFT.scala 35:12]
  assign _GEN_1017 = 9'h1f8 == cnt[8:0] ? $signed(-32'shc90) : $signed(_GEN_1016); // @[FFT.scala 35:12]
  assign _GEN_1018 = 9'h1f9 == cnt[8:0] ? $signed(-32'shafe) : $signed(_GEN_1017); // @[FFT.scala 35:12]
  assign _GEN_1019 = 9'h1fa == cnt[8:0] ? $signed(-32'sh96c) : $signed(_GEN_1018); // @[FFT.scala 35:12]
  assign _GEN_1020 = 9'h1fb == cnt[8:0] ? $signed(-32'sh7da) : $signed(_GEN_1019); // @[FFT.scala 35:12]
  assign _GEN_1021 = 9'h1fc == cnt[8:0] ? $signed(-32'sh648) : $signed(_GEN_1020); // @[FFT.scala 35:12]
  assign _GEN_1022 = 9'h1fd == cnt[8:0] ? $signed(-32'sh4b6) : $signed(_GEN_1021); // @[FFT.scala 35:12]
  assign _GEN_1023 = 9'h1fe == cnt[8:0] ? $signed(-32'sh324) : $signed(_GEN_1022); // @[FFT.scala 35:12]
  assign _GEN_2562 = 8'h1 == cnt[7:0] ? $signed(32'shfffb) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_2563 = 8'h2 == cnt[7:0] ? $signed(32'shffec) : $signed(_GEN_2562); // @[FFT.scala 34:12]
  assign _GEN_2564 = 8'h3 == cnt[7:0] ? $signed(32'shffd4) : $signed(_GEN_2563); // @[FFT.scala 34:12]
  assign _GEN_2565 = 8'h4 == cnt[7:0] ? $signed(32'shffb1) : $signed(_GEN_2564); // @[FFT.scala 34:12]
  assign _GEN_2566 = 8'h5 == cnt[7:0] ? $signed(32'shff85) : $signed(_GEN_2565); // @[FFT.scala 34:12]
  assign _GEN_2567 = 8'h6 == cnt[7:0] ? $signed(32'shff4e) : $signed(_GEN_2566); // @[FFT.scala 34:12]
  assign _GEN_2568 = 8'h7 == cnt[7:0] ? $signed(32'shff0e) : $signed(_GEN_2567); // @[FFT.scala 34:12]
  assign _GEN_2569 = 8'h8 == cnt[7:0] ? $signed(32'shfec4) : $signed(_GEN_2568); // @[FFT.scala 34:12]
  assign _GEN_2570 = 8'h9 == cnt[7:0] ? $signed(32'shfe71) : $signed(_GEN_2569); // @[FFT.scala 34:12]
  assign _GEN_2571 = 8'ha == cnt[7:0] ? $signed(32'shfe13) : $signed(_GEN_2570); // @[FFT.scala 34:12]
  assign _GEN_2572 = 8'hb == cnt[7:0] ? $signed(32'shfdac) : $signed(_GEN_2571); // @[FFT.scala 34:12]
  assign _GEN_2573 = 8'hc == cnt[7:0] ? $signed(32'shfd3b) : $signed(_GEN_2572); // @[FFT.scala 34:12]
  assign _GEN_2574 = 8'hd == cnt[7:0] ? $signed(32'shfcc0) : $signed(_GEN_2573); // @[FFT.scala 34:12]
  assign _GEN_2575 = 8'he == cnt[7:0] ? $signed(32'shfc3b) : $signed(_GEN_2574); // @[FFT.scala 34:12]
  assign _GEN_2576 = 8'hf == cnt[7:0] ? $signed(32'shfbad) : $signed(_GEN_2575); // @[FFT.scala 34:12]
  assign _GEN_2577 = 8'h10 == cnt[7:0] ? $signed(32'shfb15) : $signed(_GEN_2576); // @[FFT.scala 34:12]
  assign _GEN_2578 = 8'h11 == cnt[7:0] ? $signed(32'shfa73) : $signed(_GEN_2577); // @[FFT.scala 34:12]
  assign _GEN_2579 = 8'h12 == cnt[7:0] ? $signed(32'shf9c8) : $signed(_GEN_2578); // @[FFT.scala 34:12]
  assign _GEN_2580 = 8'h13 == cnt[7:0] ? $signed(32'shf913) : $signed(_GEN_2579); // @[FFT.scala 34:12]
  assign _GEN_2581 = 8'h14 == cnt[7:0] ? $signed(32'shf854) : $signed(_GEN_2580); // @[FFT.scala 34:12]
  assign _GEN_2582 = 8'h15 == cnt[7:0] ? $signed(32'shf78c) : $signed(_GEN_2581); // @[FFT.scala 34:12]
  assign _GEN_2583 = 8'h16 == cnt[7:0] ? $signed(32'shf6ba) : $signed(_GEN_2582); // @[FFT.scala 34:12]
  assign _GEN_2584 = 8'h17 == cnt[7:0] ? $signed(32'shf5df) : $signed(_GEN_2583); // @[FFT.scala 34:12]
  assign _GEN_2585 = 8'h18 == cnt[7:0] ? $signed(32'shf4fa) : $signed(_GEN_2584); // @[FFT.scala 34:12]
  assign _GEN_2586 = 8'h19 == cnt[7:0] ? $signed(32'shf40c) : $signed(_GEN_2585); // @[FFT.scala 34:12]
  assign _GEN_2587 = 8'h1a == cnt[7:0] ? $signed(32'shf314) : $signed(_GEN_2586); // @[FFT.scala 34:12]
  assign _GEN_2588 = 8'h1b == cnt[7:0] ? $signed(32'shf213) : $signed(_GEN_2587); // @[FFT.scala 34:12]
  assign _GEN_2589 = 8'h1c == cnt[7:0] ? $signed(32'shf109) : $signed(_GEN_2588); // @[FFT.scala 34:12]
  assign _GEN_2590 = 8'h1d == cnt[7:0] ? $signed(32'sheff5) : $signed(_GEN_2589); // @[FFT.scala 34:12]
  assign _GEN_2591 = 8'h1e == cnt[7:0] ? $signed(32'sheed9) : $signed(_GEN_2590); // @[FFT.scala 34:12]
  assign _GEN_2592 = 8'h1f == cnt[7:0] ? $signed(32'shedb3) : $signed(_GEN_2591); // @[FFT.scala 34:12]
  assign _GEN_2593 = 8'h20 == cnt[7:0] ? $signed(32'shec83) : $signed(_GEN_2592); // @[FFT.scala 34:12]
  assign _GEN_2594 = 8'h21 == cnt[7:0] ? $signed(32'sheb4b) : $signed(_GEN_2593); // @[FFT.scala 34:12]
  assign _GEN_2595 = 8'h22 == cnt[7:0] ? $signed(32'shea0a) : $signed(_GEN_2594); // @[FFT.scala 34:12]
  assign _GEN_2596 = 8'h23 == cnt[7:0] ? $signed(32'she8bf) : $signed(_GEN_2595); // @[FFT.scala 34:12]
  assign _GEN_2597 = 8'h24 == cnt[7:0] ? $signed(32'she76c) : $signed(_GEN_2596); // @[FFT.scala 34:12]
  assign _GEN_2598 = 8'h25 == cnt[7:0] ? $signed(32'she610) : $signed(_GEN_2597); // @[FFT.scala 34:12]
  assign _GEN_2599 = 8'h26 == cnt[7:0] ? $signed(32'she4aa) : $signed(_GEN_2598); // @[FFT.scala 34:12]
  assign _GEN_2600 = 8'h27 == cnt[7:0] ? $signed(32'she33c) : $signed(_GEN_2599); // @[FFT.scala 34:12]
  assign _GEN_2601 = 8'h28 == cnt[7:0] ? $signed(32'she1c6) : $signed(_GEN_2600); // @[FFT.scala 34:12]
  assign _GEN_2602 = 8'h29 == cnt[7:0] ? $signed(32'she046) : $signed(_GEN_2601); // @[FFT.scala 34:12]
  assign _GEN_2603 = 8'h2a == cnt[7:0] ? $signed(32'shdebe) : $signed(_GEN_2602); // @[FFT.scala 34:12]
  assign _GEN_2604 = 8'h2b == cnt[7:0] ? $signed(32'shdd2d) : $signed(_GEN_2603); // @[FFT.scala 34:12]
  assign _GEN_2605 = 8'h2c == cnt[7:0] ? $signed(32'shdb94) : $signed(_GEN_2604); // @[FFT.scala 34:12]
  assign _GEN_2606 = 8'h2d == cnt[7:0] ? $signed(32'shd9f2) : $signed(_GEN_2605); // @[FFT.scala 34:12]
  assign _GEN_2607 = 8'h2e == cnt[7:0] ? $signed(32'shd848) : $signed(_GEN_2606); // @[FFT.scala 34:12]
  assign _GEN_2608 = 8'h2f == cnt[7:0] ? $signed(32'shd696) : $signed(_GEN_2607); // @[FFT.scala 34:12]
  assign _GEN_2609 = 8'h30 == cnt[7:0] ? $signed(32'shd4db) : $signed(_GEN_2608); // @[FFT.scala 34:12]
  assign _GEN_2610 = 8'h31 == cnt[7:0] ? $signed(32'shd318) : $signed(_GEN_2609); // @[FFT.scala 34:12]
  assign _GEN_2611 = 8'h32 == cnt[7:0] ? $signed(32'shd14d) : $signed(_GEN_2610); // @[FFT.scala 34:12]
  assign _GEN_2612 = 8'h33 == cnt[7:0] ? $signed(32'shcf7a) : $signed(_GEN_2611); // @[FFT.scala 34:12]
  assign _GEN_2613 = 8'h34 == cnt[7:0] ? $signed(32'shcd9f) : $signed(_GEN_2612); // @[FFT.scala 34:12]
  assign _GEN_2614 = 8'h35 == cnt[7:0] ? $signed(32'shcbbc) : $signed(_GEN_2613); // @[FFT.scala 34:12]
  assign _GEN_2615 = 8'h36 == cnt[7:0] ? $signed(32'shc9d1) : $signed(_GEN_2614); // @[FFT.scala 34:12]
  assign _GEN_2616 = 8'h37 == cnt[7:0] ? $signed(32'shc7de) : $signed(_GEN_2615); // @[FFT.scala 34:12]
  assign _GEN_2617 = 8'h38 == cnt[7:0] ? $signed(32'shc5e4) : $signed(_GEN_2616); // @[FFT.scala 34:12]
  assign _GEN_2618 = 8'h39 == cnt[7:0] ? $signed(32'shc3e2) : $signed(_GEN_2617); // @[FFT.scala 34:12]
  assign _GEN_2619 = 8'h3a == cnt[7:0] ? $signed(32'shc1d8) : $signed(_GEN_2618); // @[FFT.scala 34:12]
  assign _GEN_2620 = 8'h3b == cnt[7:0] ? $signed(32'shbfc7) : $signed(_GEN_2619); // @[FFT.scala 34:12]
  assign _GEN_2621 = 8'h3c == cnt[7:0] ? $signed(32'shbdaf) : $signed(_GEN_2620); // @[FFT.scala 34:12]
  assign _GEN_2622 = 8'h3d == cnt[7:0] ? $signed(32'shbb8f) : $signed(_GEN_2621); // @[FFT.scala 34:12]
  assign _GEN_2623 = 8'h3e == cnt[7:0] ? $signed(32'shb968) : $signed(_GEN_2622); // @[FFT.scala 34:12]
  assign _GEN_2624 = 8'h3f == cnt[7:0] ? $signed(32'shb73a) : $signed(_GEN_2623); // @[FFT.scala 34:12]
  assign _GEN_2625 = 8'h40 == cnt[7:0] ? $signed(32'shb505) : $signed(_GEN_2624); // @[FFT.scala 34:12]
  assign _GEN_2626 = 8'h41 == cnt[7:0] ? $signed(32'shb2c9) : $signed(_GEN_2625); // @[FFT.scala 34:12]
  assign _GEN_2627 = 8'h42 == cnt[7:0] ? $signed(32'shb086) : $signed(_GEN_2626); // @[FFT.scala 34:12]
  assign _GEN_2628 = 8'h43 == cnt[7:0] ? $signed(32'shae3c) : $signed(_GEN_2627); // @[FFT.scala 34:12]
  assign _GEN_2629 = 8'h44 == cnt[7:0] ? $signed(32'shabeb) : $signed(_GEN_2628); // @[FFT.scala 34:12]
  assign _GEN_2630 = 8'h45 == cnt[7:0] ? $signed(32'sha994) : $signed(_GEN_2629); // @[FFT.scala 34:12]
  assign _GEN_2631 = 8'h46 == cnt[7:0] ? $signed(32'sha736) : $signed(_GEN_2630); // @[FFT.scala 34:12]
  assign _GEN_2632 = 8'h47 == cnt[7:0] ? $signed(32'sha4d2) : $signed(_GEN_2631); // @[FFT.scala 34:12]
  assign _GEN_2633 = 8'h48 == cnt[7:0] ? $signed(32'sha268) : $signed(_GEN_2632); // @[FFT.scala 34:12]
  assign _GEN_2634 = 8'h49 == cnt[7:0] ? $signed(32'sh9ff7) : $signed(_GEN_2633); // @[FFT.scala 34:12]
  assign _GEN_2635 = 8'h4a == cnt[7:0] ? $signed(32'sh9d80) : $signed(_GEN_2634); // @[FFT.scala 34:12]
  assign _GEN_2636 = 8'h4b == cnt[7:0] ? $signed(32'sh9b03) : $signed(_GEN_2635); // @[FFT.scala 34:12]
  assign _GEN_2637 = 8'h4c == cnt[7:0] ? $signed(32'sh9880) : $signed(_GEN_2636); // @[FFT.scala 34:12]
  assign _GEN_2638 = 8'h4d == cnt[7:0] ? $signed(32'sh95f7) : $signed(_GEN_2637); // @[FFT.scala 34:12]
  assign _GEN_2639 = 8'h4e == cnt[7:0] ? $signed(32'sh9368) : $signed(_GEN_2638); // @[FFT.scala 34:12]
  assign _GEN_2640 = 8'h4f == cnt[7:0] ? $signed(32'sh90d4) : $signed(_GEN_2639); // @[FFT.scala 34:12]
  assign _GEN_2641 = 8'h50 == cnt[7:0] ? $signed(32'sh8e3a) : $signed(_GEN_2640); // @[FFT.scala 34:12]
  assign _GEN_2642 = 8'h51 == cnt[7:0] ? $signed(32'sh8b9a) : $signed(_GEN_2641); // @[FFT.scala 34:12]
  assign _GEN_2643 = 8'h52 == cnt[7:0] ? $signed(32'sh88f6) : $signed(_GEN_2642); // @[FFT.scala 34:12]
  assign _GEN_2644 = 8'h53 == cnt[7:0] ? $signed(32'sh864c) : $signed(_GEN_2643); // @[FFT.scala 34:12]
  assign _GEN_2645 = 8'h54 == cnt[7:0] ? $signed(32'sh839c) : $signed(_GEN_2644); // @[FFT.scala 34:12]
  assign _GEN_2646 = 8'h55 == cnt[7:0] ? $signed(32'sh80e8) : $signed(_GEN_2645); // @[FFT.scala 34:12]
  assign _GEN_2647 = 8'h56 == cnt[7:0] ? $signed(32'sh7e2f) : $signed(_GEN_2646); // @[FFT.scala 34:12]
  assign _GEN_2648 = 8'h57 == cnt[7:0] ? $signed(32'sh7b70) : $signed(_GEN_2647); // @[FFT.scala 34:12]
  assign _GEN_2649 = 8'h58 == cnt[7:0] ? $signed(32'sh78ad) : $signed(_GEN_2648); // @[FFT.scala 34:12]
  assign _GEN_2650 = 8'h59 == cnt[7:0] ? $signed(32'sh75e6) : $signed(_GEN_2649); // @[FFT.scala 34:12]
  assign _GEN_2651 = 8'h5a == cnt[7:0] ? $signed(32'sh731a) : $signed(_GEN_2650); // @[FFT.scala 34:12]
  assign _GEN_2652 = 8'h5b == cnt[7:0] ? $signed(32'sh7049) : $signed(_GEN_2651); // @[FFT.scala 34:12]
  assign _GEN_2653 = 8'h5c == cnt[7:0] ? $signed(32'sh6d74) : $signed(_GEN_2652); // @[FFT.scala 34:12]
  assign _GEN_2654 = 8'h5d == cnt[7:0] ? $signed(32'sh6a9b) : $signed(_GEN_2653); // @[FFT.scala 34:12]
  assign _GEN_2655 = 8'h5e == cnt[7:0] ? $signed(32'sh67be) : $signed(_GEN_2654); // @[FFT.scala 34:12]
  assign _GEN_2656 = 8'h5f == cnt[7:0] ? $signed(32'sh64dd) : $signed(_GEN_2655); // @[FFT.scala 34:12]
  assign _GEN_2657 = 8'h60 == cnt[7:0] ? $signed(32'sh61f8) : $signed(_GEN_2656); // @[FFT.scala 34:12]
  assign _GEN_2658 = 8'h61 == cnt[7:0] ? $signed(32'sh5f0f) : $signed(_GEN_2657); // @[FFT.scala 34:12]
  assign _GEN_2659 = 8'h62 == cnt[7:0] ? $signed(32'sh5c22) : $signed(_GEN_2658); // @[FFT.scala 34:12]
  assign _GEN_2660 = 8'h63 == cnt[7:0] ? $signed(32'sh5932) : $signed(_GEN_2659); // @[FFT.scala 34:12]
  assign _GEN_2661 = 8'h64 == cnt[7:0] ? $signed(32'sh563e) : $signed(_GEN_2660); // @[FFT.scala 34:12]
  assign _GEN_2662 = 8'h65 == cnt[7:0] ? $signed(32'sh5348) : $signed(_GEN_2661); // @[FFT.scala 34:12]
  assign _GEN_2663 = 8'h66 == cnt[7:0] ? $signed(32'sh504d) : $signed(_GEN_2662); // @[FFT.scala 34:12]
  assign _GEN_2664 = 8'h67 == cnt[7:0] ? $signed(32'sh4d50) : $signed(_GEN_2663); // @[FFT.scala 34:12]
  assign _GEN_2665 = 8'h68 == cnt[7:0] ? $signed(32'sh4a50) : $signed(_GEN_2664); // @[FFT.scala 34:12]
  assign _GEN_2666 = 8'h69 == cnt[7:0] ? $signed(32'sh474d) : $signed(_GEN_2665); // @[FFT.scala 34:12]
  assign _GEN_2667 = 8'h6a == cnt[7:0] ? $signed(32'sh4447) : $signed(_GEN_2666); // @[FFT.scala 34:12]
  assign _GEN_2668 = 8'h6b == cnt[7:0] ? $signed(32'sh413f) : $signed(_GEN_2667); // @[FFT.scala 34:12]
  assign _GEN_2669 = 8'h6c == cnt[7:0] ? $signed(32'sh3e34) : $signed(_GEN_2668); // @[FFT.scala 34:12]
  assign _GEN_2670 = 8'h6d == cnt[7:0] ? $signed(32'sh3b27) : $signed(_GEN_2669); // @[FFT.scala 34:12]
  assign _GEN_2671 = 8'h6e == cnt[7:0] ? $signed(32'sh3817) : $signed(_GEN_2670); // @[FFT.scala 34:12]
  assign _GEN_2672 = 8'h6f == cnt[7:0] ? $signed(32'sh3505) : $signed(_GEN_2671); // @[FFT.scala 34:12]
  assign _GEN_2673 = 8'h70 == cnt[7:0] ? $signed(32'sh31f1) : $signed(_GEN_2672); // @[FFT.scala 34:12]
  assign _GEN_2674 = 8'h71 == cnt[7:0] ? $signed(32'sh2edc) : $signed(_GEN_2673); // @[FFT.scala 34:12]
  assign _GEN_2675 = 8'h72 == cnt[7:0] ? $signed(32'sh2bc4) : $signed(_GEN_2674); // @[FFT.scala 34:12]
  assign _GEN_2676 = 8'h73 == cnt[7:0] ? $signed(32'sh28ab) : $signed(_GEN_2675); // @[FFT.scala 34:12]
  assign _GEN_2677 = 8'h74 == cnt[7:0] ? $signed(32'sh2590) : $signed(_GEN_2676); // @[FFT.scala 34:12]
  assign _GEN_2678 = 8'h75 == cnt[7:0] ? $signed(32'sh2274) : $signed(_GEN_2677); // @[FFT.scala 34:12]
  assign _GEN_2679 = 8'h76 == cnt[7:0] ? $signed(32'sh1f56) : $signed(_GEN_2678); // @[FFT.scala 34:12]
  assign _GEN_2680 = 8'h77 == cnt[7:0] ? $signed(32'sh1c38) : $signed(_GEN_2679); // @[FFT.scala 34:12]
  assign _GEN_2681 = 8'h78 == cnt[7:0] ? $signed(32'sh1918) : $signed(_GEN_2680); // @[FFT.scala 34:12]
  assign _GEN_2682 = 8'h79 == cnt[7:0] ? $signed(32'sh15f7) : $signed(_GEN_2681); // @[FFT.scala 34:12]
  assign _GEN_2683 = 8'h7a == cnt[7:0] ? $signed(32'sh12d5) : $signed(_GEN_2682); // @[FFT.scala 34:12]
  assign _GEN_2684 = 8'h7b == cnt[7:0] ? $signed(32'shfb3) : $signed(_GEN_2683); // @[FFT.scala 34:12]
  assign _GEN_2685 = 8'h7c == cnt[7:0] ? $signed(32'shc90) : $signed(_GEN_2684); // @[FFT.scala 34:12]
  assign _GEN_2686 = 8'h7d == cnt[7:0] ? $signed(32'sh96c) : $signed(_GEN_2685); // @[FFT.scala 34:12]
  assign _GEN_2687 = 8'h7e == cnt[7:0] ? $signed(32'sh648) : $signed(_GEN_2686); // @[FFT.scala 34:12]
  assign _GEN_2688 = 8'h7f == cnt[7:0] ? $signed(32'sh324) : $signed(_GEN_2687); // @[FFT.scala 34:12]
  assign _GEN_2689 = 8'h80 == cnt[7:0] ? $signed(32'sh0) : $signed(_GEN_2688); // @[FFT.scala 34:12]
  assign _GEN_2690 = 8'h81 == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_2689); // @[FFT.scala 34:12]
  assign _GEN_2691 = 8'h82 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_2690); // @[FFT.scala 34:12]
  assign _GEN_2692 = 8'h83 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_2691); // @[FFT.scala 34:12]
  assign _GEN_2693 = 8'h84 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_2692); // @[FFT.scala 34:12]
  assign _GEN_2694 = 8'h85 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_2693); // @[FFT.scala 34:12]
  assign _GEN_2695 = 8'h86 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_2694); // @[FFT.scala 34:12]
  assign _GEN_2696 = 8'h87 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_2695); // @[FFT.scala 34:12]
  assign _GEN_2697 = 8'h88 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_2696); // @[FFT.scala 34:12]
  assign _GEN_2698 = 8'h89 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_2697); // @[FFT.scala 34:12]
  assign _GEN_2699 = 8'h8a == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_2698); // @[FFT.scala 34:12]
  assign _GEN_2700 = 8'h8b == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_2699); // @[FFT.scala 34:12]
  assign _GEN_2701 = 8'h8c == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_2700); // @[FFT.scala 34:12]
  assign _GEN_2702 = 8'h8d == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_2701); // @[FFT.scala 34:12]
  assign _GEN_2703 = 8'h8e == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2702); // @[FFT.scala 34:12]
  assign _GEN_2704 = 8'h8f == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_2703); // @[FFT.scala 34:12]
  assign _GEN_2705 = 8'h90 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_2704); // @[FFT.scala 34:12]
  assign _GEN_2706 = 8'h91 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_2705); // @[FFT.scala 34:12]
  assign _GEN_2707 = 8'h92 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_2706); // @[FFT.scala 34:12]
  assign _GEN_2708 = 8'h93 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_2707); // @[FFT.scala 34:12]
  assign _GEN_2709 = 8'h94 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_2708); // @[FFT.scala 34:12]
  assign _GEN_2710 = 8'h95 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_2709); // @[FFT.scala 34:12]
  assign _GEN_2711 = 8'h96 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_2710); // @[FFT.scala 34:12]
  assign _GEN_2712 = 8'h97 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_2711); // @[FFT.scala 34:12]
  assign _GEN_2713 = 8'h98 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_2712); // @[FFT.scala 34:12]
  assign _GEN_2714 = 8'h99 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_2713); // @[FFT.scala 34:12]
  assign _GEN_2715 = 8'h9a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_2714); // @[FFT.scala 34:12]
  assign _GEN_2716 = 8'h9b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_2715); // @[FFT.scala 34:12]
  assign _GEN_2717 = 8'h9c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_2716); // @[FFT.scala 34:12]
  assign _GEN_2718 = 8'h9d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_2717); // @[FFT.scala 34:12]
  assign _GEN_2719 = 8'h9e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_2718); // @[FFT.scala 34:12]
  assign _GEN_2720 = 8'h9f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_2719); // @[FFT.scala 34:12]
  assign _GEN_2721 = 8'ha0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_2720); // @[FFT.scala 34:12]
  assign _GEN_2722 = 8'ha1 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_2721); // @[FFT.scala 34:12]
  assign _GEN_2723 = 8'ha2 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_2722); // @[FFT.scala 34:12]
  assign _GEN_2724 = 8'ha3 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_2723); // @[FFT.scala 34:12]
  assign _GEN_2725 = 8'ha4 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_2724); // @[FFT.scala 34:12]
  assign _GEN_2726 = 8'ha5 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_2725); // @[FFT.scala 34:12]
  assign _GEN_2727 = 8'ha6 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_2726); // @[FFT.scala 34:12]
  assign _GEN_2728 = 8'ha7 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_2727); // @[FFT.scala 34:12]
  assign _GEN_2729 = 8'ha8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_2728); // @[FFT.scala 34:12]
  assign _GEN_2730 = 8'ha9 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_2729); // @[FFT.scala 34:12]
  assign _GEN_2731 = 8'haa == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2730); // @[FFT.scala 34:12]
  assign _GEN_2732 = 8'hab == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_2731); // @[FFT.scala 34:12]
  assign _GEN_2733 = 8'hac == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_2732); // @[FFT.scala 34:12]
  assign _GEN_2734 = 8'had == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_2733); // @[FFT.scala 34:12]
  assign _GEN_2735 = 8'hae == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_2734); // @[FFT.scala 34:12]
  assign _GEN_2736 = 8'haf == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_2735); // @[FFT.scala 34:12]
  assign _GEN_2737 = 8'hb0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2736); // @[FFT.scala 34:12]
  assign _GEN_2738 = 8'hb1 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_2737); // @[FFT.scala 34:12]
  assign _GEN_2739 = 8'hb2 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_2738); // @[FFT.scala 34:12]
  assign _GEN_2740 = 8'hb3 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_2739); // @[FFT.scala 34:12]
  assign _GEN_2741 = 8'hb4 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_2740); // @[FFT.scala 34:12]
  assign _GEN_2742 = 8'hb5 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_2741); // @[FFT.scala 34:12]
  assign _GEN_2743 = 8'hb6 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_2742); // @[FFT.scala 34:12]
  assign _GEN_2744 = 8'hb7 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_2743); // @[FFT.scala 34:12]
  assign _GEN_2745 = 8'hb8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_2744); // @[FFT.scala 34:12]
  assign _GEN_2746 = 8'hb9 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_2745); // @[FFT.scala 34:12]
  assign _GEN_2747 = 8'hba == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_2746); // @[FFT.scala 34:12]
  assign _GEN_2748 = 8'hbb == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_2747); // @[FFT.scala 34:12]
  assign _GEN_2749 = 8'hbc == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_2748); // @[FFT.scala 34:12]
  assign _GEN_2750 = 8'hbd == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_2749); // @[FFT.scala 34:12]
  assign _GEN_2751 = 8'hbe == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_2750); // @[FFT.scala 34:12]
  assign _GEN_2752 = 8'hbf == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_2751); // @[FFT.scala 34:12]
  assign _GEN_2753 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_2752); // @[FFT.scala 34:12]
  assign _GEN_2754 = 8'hc1 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_2753); // @[FFT.scala 34:12]
  assign _GEN_2755 = 8'hc2 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_2754); // @[FFT.scala 34:12]
  assign _GEN_2756 = 8'hc3 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_2755); // @[FFT.scala 34:12]
  assign _GEN_2757 = 8'hc4 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_2756); // @[FFT.scala 34:12]
  assign _GEN_2758 = 8'hc5 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_2757); // @[FFT.scala 34:12]
  assign _GEN_2759 = 8'hc6 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_2758); // @[FFT.scala 34:12]
  assign _GEN_2760 = 8'hc7 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_2759); // @[FFT.scala 34:12]
  assign _GEN_2761 = 8'hc8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_2760); // @[FFT.scala 34:12]
  assign _GEN_2762 = 8'hc9 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_2761); // @[FFT.scala 34:12]
  assign _GEN_2763 = 8'hca == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_2762); // @[FFT.scala 34:12]
  assign _GEN_2764 = 8'hcb == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_2763); // @[FFT.scala 34:12]
  assign _GEN_2765 = 8'hcc == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_2764); // @[FFT.scala 34:12]
  assign _GEN_2766 = 8'hcd == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_2765); // @[FFT.scala 34:12]
  assign _GEN_2767 = 8'hce == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_2766); // @[FFT.scala 34:12]
  assign _GEN_2768 = 8'hcf == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_2767); // @[FFT.scala 34:12]
  assign _GEN_2769 = 8'hd0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_2768); // @[FFT.scala 34:12]
  assign _GEN_2770 = 8'hd1 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_2769); // @[FFT.scala 34:12]
  assign _GEN_2771 = 8'hd2 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_2770); // @[FFT.scala 34:12]
  assign _GEN_2772 = 8'hd3 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_2771); // @[FFT.scala 34:12]
  assign _GEN_2773 = 8'hd4 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_2772); // @[FFT.scala 34:12]
  assign _GEN_2774 = 8'hd5 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_2773); // @[FFT.scala 34:12]
  assign _GEN_2775 = 8'hd6 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_2774); // @[FFT.scala 34:12]
  assign _GEN_2776 = 8'hd7 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_2775); // @[FFT.scala 34:12]
  assign _GEN_2777 = 8'hd8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_2776); // @[FFT.scala 34:12]
  assign _GEN_2778 = 8'hd9 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_2777); // @[FFT.scala 34:12]
  assign _GEN_2779 = 8'hda == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_2778); // @[FFT.scala 34:12]
  assign _GEN_2780 = 8'hdb == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_2779); // @[FFT.scala 34:12]
  assign _GEN_2781 = 8'hdc == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_2780); // @[FFT.scala 34:12]
  assign _GEN_2782 = 8'hdd == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_2781); // @[FFT.scala 34:12]
  assign _GEN_2783 = 8'hde == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_2782); // @[FFT.scala 34:12]
  assign _GEN_2784 = 8'hdf == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_2783); // @[FFT.scala 34:12]
  assign _GEN_2785 = 8'he0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_2784); // @[FFT.scala 34:12]
  assign _GEN_2786 = 8'he1 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_2785); // @[FFT.scala 34:12]
  assign _GEN_2787 = 8'he2 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_2786); // @[FFT.scala 34:12]
  assign _GEN_2788 = 8'he3 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_2787); // @[FFT.scala 34:12]
  assign _GEN_2789 = 8'he4 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_2788); // @[FFT.scala 34:12]
  assign _GEN_2790 = 8'he5 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_2789); // @[FFT.scala 34:12]
  assign _GEN_2791 = 8'he6 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_2790); // @[FFT.scala 34:12]
  assign _GEN_2792 = 8'he7 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_2791); // @[FFT.scala 34:12]
  assign _GEN_2793 = 8'he8 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_2792); // @[FFT.scala 34:12]
  assign _GEN_2794 = 8'he9 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_2793); // @[FFT.scala 34:12]
  assign _GEN_2795 = 8'hea == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_2794); // @[FFT.scala 34:12]
  assign _GEN_2796 = 8'heb == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_2795); // @[FFT.scala 34:12]
  assign _GEN_2797 = 8'hec == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_2796); // @[FFT.scala 34:12]
  assign _GEN_2798 = 8'hed == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_2797); // @[FFT.scala 34:12]
  assign _GEN_2799 = 8'hee == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_2798); // @[FFT.scala 34:12]
  assign _GEN_2800 = 8'hef == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_2799); // @[FFT.scala 34:12]
  assign _GEN_2801 = 8'hf0 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_2800); // @[FFT.scala 34:12]
  assign _GEN_2802 = 8'hf1 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_2801); // @[FFT.scala 34:12]
  assign _GEN_2803 = 8'hf2 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_2802); // @[FFT.scala 34:12]
  assign _GEN_2804 = 8'hf3 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_2803); // @[FFT.scala 34:12]
  assign _GEN_2805 = 8'hf4 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_2804); // @[FFT.scala 34:12]
  assign _GEN_2806 = 8'hf5 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_2805); // @[FFT.scala 34:12]
  assign _GEN_2807 = 8'hf6 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_2806); // @[FFT.scala 34:12]
  assign _GEN_2808 = 8'hf7 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_2807); // @[FFT.scala 34:12]
  assign _GEN_2809 = 8'hf8 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_2808); // @[FFT.scala 34:12]
  assign _GEN_2810 = 8'hf9 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_2809); // @[FFT.scala 34:12]
  assign _GEN_2811 = 8'hfa == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_2810); // @[FFT.scala 34:12]
  assign _GEN_2812 = 8'hfb == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_2811); // @[FFT.scala 34:12]
  assign _GEN_2813 = 8'hfc == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_2812); // @[FFT.scala 34:12]
  assign _GEN_2814 = 8'hfd == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_2813); // @[FFT.scala 34:12]
  assign _GEN_2815 = 8'hfe == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_2814); // @[FFT.scala 34:12]
  assign _GEN_2818 = 8'h1 == cnt[7:0] ? $signed(-32'sh324) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_2819 = 8'h2 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_2818); // @[FFT.scala 35:12]
  assign _GEN_2820 = 8'h3 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_2819); // @[FFT.scala 35:12]
  assign _GEN_2821 = 8'h4 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_2820); // @[FFT.scala 35:12]
  assign _GEN_2822 = 8'h5 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_2821); // @[FFT.scala 35:12]
  assign _GEN_2823 = 8'h6 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_2822); // @[FFT.scala 35:12]
  assign _GEN_2824 = 8'h7 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_2823); // @[FFT.scala 35:12]
  assign _GEN_2825 = 8'h8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_2824); // @[FFT.scala 35:12]
  assign _GEN_2826 = 8'h9 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_2825); // @[FFT.scala 35:12]
  assign _GEN_2827 = 8'ha == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_2826); // @[FFT.scala 35:12]
  assign _GEN_2828 = 8'hb == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_2827); // @[FFT.scala 35:12]
  assign _GEN_2829 = 8'hc == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_2828); // @[FFT.scala 35:12]
  assign _GEN_2830 = 8'hd == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_2829); // @[FFT.scala 35:12]
  assign _GEN_2831 = 8'he == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2830); // @[FFT.scala 35:12]
  assign _GEN_2832 = 8'hf == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_2831); // @[FFT.scala 35:12]
  assign _GEN_2833 = 8'h10 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_2832); // @[FFT.scala 35:12]
  assign _GEN_2834 = 8'h11 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_2833); // @[FFT.scala 35:12]
  assign _GEN_2835 = 8'h12 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_2834); // @[FFT.scala 35:12]
  assign _GEN_2836 = 8'h13 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_2835); // @[FFT.scala 35:12]
  assign _GEN_2837 = 8'h14 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_2836); // @[FFT.scala 35:12]
  assign _GEN_2838 = 8'h15 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_2837); // @[FFT.scala 35:12]
  assign _GEN_2839 = 8'h16 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_2838); // @[FFT.scala 35:12]
  assign _GEN_2840 = 8'h17 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_2839); // @[FFT.scala 35:12]
  assign _GEN_2841 = 8'h18 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_2840); // @[FFT.scala 35:12]
  assign _GEN_2842 = 8'h19 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_2841); // @[FFT.scala 35:12]
  assign _GEN_2843 = 8'h1a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_2842); // @[FFT.scala 35:12]
  assign _GEN_2844 = 8'h1b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_2843); // @[FFT.scala 35:12]
  assign _GEN_2845 = 8'h1c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_2844); // @[FFT.scala 35:12]
  assign _GEN_2846 = 8'h1d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_2845); // @[FFT.scala 35:12]
  assign _GEN_2847 = 8'h1e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_2846); // @[FFT.scala 35:12]
  assign _GEN_2848 = 8'h1f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_2847); // @[FFT.scala 35:12]
  assign _GEN_2849 = 8'h20 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_2848); // @[FFT.scala 35:12]
  assign _GEN_2850 = 8'h21 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_2849); // @[FFT.scala 35:12]
  assign _GEN_2851 = 8'h22 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_2850); // @[FFT.scala 35:12]
  assign _GEN_2852 = 8'h23 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_2851); // @[FFT.scala 35:12]
  assign _GEN_2853 = 8'h24 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_2852); // @[FFT.scala 35:12]
  assign _GEN_2854 = 8'h25 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_2853); // @[FFT.scala 35:12]
  assign _GEN_2855 = 8'h26 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_2854); // @[FFT.scala 35:12]
  assign _GEN_2856 = 8'h27 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_2855); // @[FFT.scala 35:12]
  assign _GEN_2857 = 8'h28 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_2856); // @[FFT.scala 35:12]
  assign _GEN_2858 = 8'h29 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_2857); // @[FFT.scala 35:12]
  assign _GEN_2859 = 8'h2a == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2858); // @[FFT.scala 35:12]
  assign _GEN_2860 = 8'h2b == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_2859); // @[FFT.scala 35:12]
  assign _GEN_2861 = 8'h2c == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_2860); // @[FFT.scala 35:12]
  assign _GEN_2862 = 8'h2d == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_2861); // @[FFT.scala 35:12]
  assign _GEN_2863 = 8'h2e == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_2862); // @[FFT.scala 35:12]
  assign _GEN_2864 = 8'h2f == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_2863); // @[FFT.scala 35:12]
  assign _GEN_2865 = 8'h30 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2864); // @[FFT.scala 35:12]
  assign _GEN_2866 = 8'h31 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_2865); // @[FFT.scala 35:12]
  assign _GEN_2867 = 8'h32 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_2866); // @[FFT.scala 35:12]
  assign _GEN_2868 = 8'h33 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_2867); // @[FFT.scala 35:12]
  assign _GEN_2869 = 8'h34 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_2868); // @[FFT.scala 35:12]
  assign _GEN_2870 = 8'h35 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_2869); // @[FFT.scala 35:12]
  assign _GEN_2871 = 8'h36 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_2870); // @[FFT.scala 35:12]
  assign _GEN_2872 = 8'h37 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_2871); // @[FFT.scala 35:12]
  assign _GEN_2873 = 8'h38 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_2872); // @[FFT.scala 35:12]
  assign _GEN_2874 = 8'h39 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_2873); // @[FFT.scala 35:12]
  assign _GEN_2875 = 8'h3a == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_2874); // @[FFT.scala 35:12]
  assign _GEN_2876 = 8'h3b == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_2875); // @[FFT.scala 35:12]
  assign _GEN_2877 = 8'h3c == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_2876); // @[FFT.scala 35:12]
  assign _GEN_2878 = 8'h3d == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_2877); // @[FFT.scala 35:12]
  assign _GEN_2879 = 8'h3e == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_2878); // @[FFT.scala 35:12]
  assign _GEN_2880 = 8'h3f == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_2879); // @[FFT.scala 35:12]
  assign _GEN_2881 = 8'h40 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_2880); // @[FFT.scala 35:12]
  assign _GEN_2882 = 8'h41 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_2881); // @[FFT.scala 35:12]
  assign _GEN_2883 = 8'h42 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_2882); // @[FFT.scala 35:12]
  assign _GEN_2884 = 8'h43 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_2883); // @[FFT.scala 35:12]
  assign _GEN_2885 = 8'h44 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_2884); // @[FFT.scala 35:12]
  assign _GEN_2886 = 8'h45 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_2885); // @[FFT.scala 35:12]
  assign _GEN_2887 = 8'h46 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_2886); // @[FFT.scala 35:12]
  assign _GEN_2888 = 8'h47 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_2887); // @[FFT.scala 35:12]
  assign _GEN_2889 = 8'h48 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_2888); // @[FFT.scala 35:12]
  assign _GEN_2890 = 8'h49 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_2889); // @[FFT.scala 35:12]
  assign _GEN_2891 = 8'h4a == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_2890); // @[FFT.scala 35:12]
  assign _GEN_2892 = 8'h4b == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_2891); // @[FFT.scala 35:12]
  assign _GEN_2893 = 8'h4c == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_2892); // @[FFT.scala 35:12]
  assign _GEN_2894 = 8'h4d == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_2893); // @[FFT.scala 35:12]
  assign _GEN_2895 = 8'h4e == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_2894); // @[FFT.scala 35:12]
  assign _GEN_2896 = 8'h4f == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_2895); // @[FFT.scala 35:12]
  assign _GEN_2897 = 8'h50 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_2896); // @[FFT.scala 35:12]
  assign _GEN_2898 = 8'h51 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_2897); // @[FFT.scala 35:12]
  assign _GEN_2899 = 8'h52 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_2898); // @[FFT.scala 35:12]
  assign _GEN_2900 = 8'h53 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_2899); // @[FFT.scala 35:12]
  assign _GEN_2901 = 8'h54 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_2900); // @[FFT.scala 35:12]
  assign _GEN_2902 = 8'h55 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_2901); // @[FFT.scala 35:12]
  assign _GEN_2903 = 8'h56 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_2902); // @[FFT.scala 35:12]
  assign _GEN_2904 = 8'h57 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_2903); // @[FFT.scala 35:12]
  assign _GEN_2905 = 8'h58 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_2904); // @[FFT.scala 35:12]
  assign _GEN_2906 = 8'h59 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_2905); // @[FFT.scala 35:12]
  assign _GEN_2907 = 8'h5a == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_2906); // @[FFT.scala 35:12]
  assign _GEN_2908 = 8'h5b == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_2907); // @[FFT.scala 35:12]
  assign _GEN_2909 = 8'h5c == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_2908); // @[FFT.scala 35:12]
  assign _GEN_2910 = 8'h5d == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_2909); // @[FFT.scala 35:12]
  assign _GEN_2911 = 8'h5e == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_2910); // @[FFT.scala 35:12]
  assign _GEN_2912 = 8'h5f == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_2911); // @[FFT.scala 35:12]
  assign _GEN_2913 = 8'h60 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_2912); // @[FFT.scala 35:12]
  assign _GEN_2914 = 8'h61 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_2913); // @[FFT.scala 35:12]
  assign _GEN_2915 = 8'h62 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_2914); // @[FFT.scala 35:12]
  assign _GEN_2916 = 8'h63 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_2915); // @[FFT.scala 35:12]
  assign _GEN_2917 = 8'h64 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_2916); // @[FFT.scala 35:12]
  assign _GEN_2918 = 8'h65 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_2917); // @[FFT.scala 35:12]
  assign _GEN_2919 = 8'h66 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_2918); // @[FFT.scala 35:12]
  assign _GEN_2920 = 8'h67 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_2919); // @[FFT.scala 35:12]
  assign _GEN_2921 = 8'h68 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_2920); // @[FFT.scala 35:12]
  assign _GEN_2922 = 8'h69 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_2921); // @[FFT.scala 35:12]
  assign _GEN_2923 = 8'h6a == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_2922); // @[FFT.scala 35:12]
  assign _GEN_2924 = 8'h6b == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_2923); // @[FFT.scala 35:12]
  assign _GEN_2925 = 8'h6c == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_2924); // @[FFT.scala 35:12]
  assign _GEN_2926 = 8'h6d == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_2925); // @[FFT.scala 35:12]
  assign _GEN_2927 = 8'h6e == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_2926); // @[FFT.scala 35:12]
  assign _GEN_2928 = 8'h6f == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_2927); // @[FFT.scala 35:12]
  assign _GEN_2929 = 8'h70 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_2928); // @[FFT.scala 35:12]
  assign _GEN_2930 = 8'h71 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_2929); // @[FFT.scala 35:12]
  assign _GEN_2931 = 8'h72 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_2930); // @[FFT.scala 35:12]
  assign _GEN_2932 = 8'h73 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_2931); // @[FFT.scala 35:12]
  assign _GEN_2933 = 8'h74 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_2932); // @[FFT.scala 35:12]
  assign _GEN_2934 = 8'h75 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_2933); // @[FFT.scala 35:12]
  assign _GEN_2935 = 8'h76 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_2934); // @[FFT.scala 35:12]
  assign _GEN_2936 = 8'h77 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_2935); // @[FFT.scala 35:12]
  assign _GEN_2937 = 8'h78 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_2936); // @[FFT.scala 35:12]
  assign _GEN_2938 = 8'h79 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_2937); // @[FFT.scala 35:12]
  assign _GEN_2939 = 8'h7a == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_2938); // @[FFT.scala 35:12]
  assign _GEN_2940 = 8'h7b == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_2939); // @[FFT.scala 35:12]
  assign _GEN_2941 = 8'h7c == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_2940); // @[FFT.scala 35:12]
  assign _GEN_2942 = 8'h7d == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_2941); // @[FFT.scala 35:12]
  assign _GEN_2943 = 8'h7e == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_2942); // @[FFT.scala 35:12]
  assign _GEN_2944 = 8'h7f == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_2943); // @[FFT.scala 35:12]
  assign _GEN_2945 = 8'h80 == cnt[7:0] ? $signed(-32'sh10000) : $signed(_GEN_2944); // @[FFT.scala 35:12]
  assign _GEN_2946 = 8'h81 == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_2945); // @[FFT.scala 35:12]
  assign _GEN_2947 = 8'h82 == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_2946); // @[FFT.scala 35:12]
  assign _GEN_2948 = 8'h83 == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_2947); // @[FFT.scala 35:12]
  assign _GEN_2949 = 8'h84 == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_2948); // @[FFT.scala 35:12]
  assign _GEN_2950 = 8'h85 == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_2949); // @[FFT.scala 35:12]
  assign _GEN_2951 = 8'h86 == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_2950); // @[FFT.scala 35:12]
  assign _GEN_2952 = 8'h87 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_2951); // @[FFT.scala 35:12]
  assign _GEN_2953 = 8'h88 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_2952); // @[FFT.scala 35:12]
  assign _GEN_2954 = 8'h89 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_2953); // @[FFT.scala 35:12]
  assign _GEN_2955 = 8'h8a == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_2954); // @[FFT.scala 35:12]
  assign _GEN_2956 = 8'h8b == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_2955); // @[FFT.scala 35:12]
  assign _GEN_2957 = 8'h8c == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_2956); // @[FFT.scala 35:12]
  assign _GEN_2958 = 8'h8d == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_2957); // @[FFT.scala 35:12]
  assign _GEN_2959 = 8'h8e == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_2958); // @[FFT.scala 35:12]
  assign _GEN_2960 = 8'h8f == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_2959); // @[FFT.scala 35:12]
  assign _GEN_2961 = 8'h90 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_2960); // @[FFT.scala 35:12]
  assign _GEN_2962 = 8'h91 == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_2961); // @[FFT.scala 35:12]
  assign _GEN_2963 = 8'h92 == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_2962); // @[FFT.scala 35:12]
  assign _GEN_2964 = 8'h93 == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_2963); // @[FFT.scala 35:12]
  assign _GEN_2965 = 8'h94 == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_2964); // @[FFT.scala 35:12]
  assign _GEN_2966 = 8'h95 == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_2965); // @[FFT.scala 35:12]
  assign _GEN_2967 = 8'h96 == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_2966); // @[FFT.scala 35:12]
  assign _GEN_2968 = 8'h97 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_2967); // @[FFT.scala 35:12]
  assign _GEN_2969 = 8'h98 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_2968); // @[FFT.scala 35:12]
  assign _GEN_2970 = 8'h99 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_2969); // @[FFT.scala 35:12]
  assign _GEN_2971 = 8'h9a == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_2970); // @[FFT.scala 35:12]
  assign _GEN_2972 = 8'h9b == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_2971); // @[FFT.scala 35:12]
  assign _GEN_2973 = 8'h9c == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_2972); // @[FFT.scala 35:12]
  assign _GEN_2974 = 8'h9d == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_2973); // @[FFT.scala 35:12]
  assign _GEN_2975 = 8'h9e == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_2974); // @[FFT.scala 35:12]
  assign _GEN_2976 = 8'h9f == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_2975); // @[FFT.scala 35:12]
  assign _GEN_2977 = 8'ha0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_2976); // @[FFT.scala 35:12]
  assign _GEN_2978 = 8'ha1 == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_2977); // @[FFT.scala 35:12]
  assign _GEN_2979 = 8'ha2 == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_2978); // @[FFT.scala 35:12]
  assign _GEN_2980 = 8'ha3 == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_2979); // @[FFT.scala 35:12]
  assign _GEN_2981 = 8'ha4 == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_2980); // @[FFT.scala 35:12]
  assign _GEN_2982 = 8'ha5 == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_2981); // @[FFT.scala 35:12]
  assign _GEN_2983 = 8'ha6 == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_2982); // @[FFT.scala 35:12]
  assign _GEN_2984 = 8'ha7 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_2983); // @[FFT.scala 35:12]
  assign _GEN_2985 = 8'ha8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_2984); // @[FFT.scala 35:12]
  assign _GEN_2986 = 8'ha9 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_2985); // @[FFT.scala 35:12]
  assign _GEN_2987 = 8'haa == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_2986); // @[FFT.scala 35:12]
  assign _GEN_2988 = 8'hab == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_2987); // @[FFT.scala 35:12]
  assign _GEN_2989 = 8'hac == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_2988); // @[FFT.scala 35:12]
  assign _GEN_2990 = 8'had == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_2989); // @[FFT.scala 35:12]
  assign _GEN_2991 = 8'hae == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_2990); // @[FFT.scala 35:12]
  assign _GEN_2992 = 8'haf == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_2991); // @[FFT.scala 35:12]
  assign _GEN_2993 = 8'hb0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_2992); // @[FFT.scala 35:12]
  assign _GEN_2994 = 8'hb1 == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_2993); // @[FFT.scala 35:12]
  assign _GEN_2995 = 8'hb2 == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_2994); // @[FFT.scala 35:12]
  assign _GEN_2996 = 8'hb3 == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_2995); // @[FFT.scala 35:12]
  assign _GEN_2997 = 8'hb4 == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_2996); // @[FFT.scala 35:12]
  assign _GEN_2998 = 8'hb5 == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_2997); // @[FFT.scala 35:12]
  assign _GEN_2999 = 8'hb6 == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_2998); // @[FFT.scala 35:12]
  assign _GEN_3000 = 8'hb7 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_2999); // @[FFT.scala 35:12]
  assign _GEN_3001 = 8'hb8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_3000); // @[FFT.scala 35:12]
  assign _GEN_3002 = 8'hb9 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_3001); // @[FFT.scala 35:12]
  assign _GEN_3003 = 8'hba == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_3002); // @[FFT.scala 35:12]
  assign _GEN_3004 = 8'hbb == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_3003); // @[FFT.scala 35:12]
  assign _GEN_3005 = 8'hbc == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_3004); // @[FFT.scala 35:12]
  assign _GEN_3006 = 8'hbd == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_3005); // @[FFT.scala 35:12]
  assign _GEN_3007 = 8'hbe == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_3006); // @[FFT.scala 35:12]
  assign _GEN_3008 = 8'hbf == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_3007); // @[FFT.scala 35:12]
  assign _GEN_3009 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_3008); // @[FFT.scala 35:12]
  assign _GEN_3010 = 8'hc1 == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_3009); // @[FFT.scala 35:12]
  assign _GEN_3011 = 8'hc2 == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_3010); // @[FFT.scala 35:12]
  assign _GEN_3012 = 8'hc3 == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_3011); // @[FFT.scala 35:12]
  assign _GEN_3013 = 8'hc4 == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_3012); // @[FFT.scala 35:12]
  assign _GEN_3014 = 8'hc5 == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_3013); // @[FFT.scala 35:12]
  assign _GEN_3015 = 8'hc6 == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_3014); // @[FFT.scala 35:12]
  assign _GEN_3016 = 8'hc7 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_3015); // @[FFT.scala 35:12]
  assign _GEN_3017 = 8'hc8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_3016); // @[FFT.scala 35:12]
  assign _GEN_3018 = 8'hc9 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_3017); // @[FFT.scala 35:12]
  assign _GEN_3019 = 8'hca == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_3018); // @[FFT.scala 35:12]
  assign _GEN_3020 = 8'hcb == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_3019); // @[FFT.scala 35:12]
  assign _GEN_3021 = 8'hcc == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_3020); // @[FFT.scala 35:12]
  assign _GEN_3022 = 8'hcd == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_3021); // @[FFT.scala 35:12]
  assign _GEN_3023 = 8'hce == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_3022); // @[FFT.scala 35:12]
  assign _GEN_3024 = 8'hcf == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_3023); // @[FFT.scala 35:12]
  assign _GEN_3025 = 8'hd0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3024); // @[FFT.scala 35:12]
  assign _GEN_3026 = 8'hd1 == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_3025); // @[FFT.scala 35:12]
  assign _GEN_3027 = 8'hd2 == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_3026); // @[FFT.scala 35:12]
  assign _GEN_3028 = 8'hd3 == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_3027); // @[FFT.scala 35:12]
  assign _GEN_3029 = 8'hd4 == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_3028); // @[FFT.scala 35:12]
  assign _GEN_3030 = 8'hd5 == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_3029); // @[FFT.scala 35:12]
  assign _GEN_3031 = 8'hd6 == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_3030); // @[FFT.scala 35:12]
  assign _GEN_3032 = 8'hd7 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_3031); // @[FFT.scala 35:12]
  assign _GEN_3033 = 8'hd8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_3032); // @[FFT.scala 35:12]
  assign _GEN_3034 = 8'hd9 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_3033); // @[FFT.scala 35:12]
  assign _GEN_3035 = 8'hda == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_3034); // @[FFT.scala 35:12]
  assign _GEN_3036 = 8'hdb == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_3035); // @[FFT.scala 35:12]
  assign _GEN_3037 = 8'hdc == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_3036); // @[FFT.scala 35:12]
  assign _GEN_3038 = 8'hdd == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_3037); // @[FFT.scala 35:12]
  assign _GEN_3039 = 8'hde == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_3038); // @[FFT.scala 35:12]
  assign _GEN_3040 = 8'hdf == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_3039); // @[FFT.scala 35:12]
  assign _GEN_3041 = 8'he0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_3040); // @[FFT.scala 35:12]
  assign _GEN_3042 = 8'he1 == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_3041); // @[FFT.scala 35:12]
  assign _GEN_3043 = 8'he2 == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_3042); // @[FFT.scala 35:12]
  assign _GEN_3044 = 8'he3 == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_3043); // @[FFT.scala 35:12]
  assign _GEN_3045 = 8'he4 == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_3044); // @[FFT.scala 35:12]
  assign _GEN_3046 = 8'he5 == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_3045); // @[FFT.scala 35:12]
  assign _GEN_3047 = 8'he6 == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_3046); // @[FFT.scala 35:12]
  assign _GEN_3048 = 8'he7 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_3047); // @[FFT.scala 35:12]
  assign _GEN_3049 = 8'he8 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_3048); // @[FFT.scala 35:12]
  assign _GEN_3050 = 8'he9 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_3049); // @[FFT.scala 35:12]
  assign _GEN_3051 = 8'hea == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_3050); // @[FFT.scala 35:12]
  assign _GEN_3052 = 8'heb == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_3051); // @[FFT.scala 35:12]
  assign _GEN_3053 = 8'hec == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_3052); // @[FFT.scala 35:12]
  assign _GEN_3054 = 8'hed == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_3053); // @[FFT.scala 35:12]
  assign _GEN_3055 = 8'hee == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_3054); // @[FFT.scala 35:12]
  assign _GEN_3056 = 8'hef == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_3055); // @[FFT.scala 35:12]
  assign _GEN_3057 = 8'hf0 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_3056); // @[FFT.scala 35:12]
  assign _GEN_3058 = 8'hf1 == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_3057); // @[FFT.scala 35:12]
  assign _GEN_3059 = 8'hf2 == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_3058); // @[FFT.scala 35:12]
  assign _GEN_3060 = 8'hf3 == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_3059); // @[FFT.scala 35:12]
  assign _GEN_3061 = 8'hf4 == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_3060); // @[FFT.scala 35:12]
  assign _GEN_3062 = 8'hf5 == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_3061); // @[FFT.scala 35:12]
  assign _GEN_3063 = 8'hf6 == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_3062); // @[FFT.scala 35:12]
  assign _GEN_3064 = 8'hf7 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_3063); // @[FFT.scala 35:12]
  assign _GEN_3065 = 8'hf8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_3064); // @[FFT.scala 35:12]
  assign _GEN_3066 = 8'hf9 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_3065); // @[FFT.scala 35:12]
  assign _GEN_3067 = 8'hfa == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_3066); // @[FFT.scala 35:12]
  assign _GEN_3068 = 8'hfb == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_3067); // @[FFT.scala 35:12]
  assign _GEN_3069 = 8'hfc == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_3068); // @[FFT.scala 35:12]
  assign _GEN_3070 = 8'hfd == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_3069); // @[FFT.scala 35:12]
  assign _GEN_3071 = 8'hfe == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_3070); // @[FFT.scala 35:12]
  assign _GEN_3842 = 7'h1 == cnt[6:0] ? $signed(32'shffec) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_3843 = 7'h2 == cnt[6:0] ? $signed(32'shffb1) : $signed(_GEN_3842); // @[FFT.scala 34:12]
  assign _GEN_3844 = 7'h3 == cnt[6:0] ? $signed(32'shff4e) : $signed(_GEN_3843); // @[FFT.scala 34:12]
  assign _GEN_3845 = 7'h4 == cnt[6:0] ? $signed(32'shfec4) : $signed(_GEN_3844); // @[FFT.scala 34:12]
  assign _GEN_3846 = 7'h5 == cnt[6:0] ? $signed(32'shfe13) : $signed(_GEN_3845); // @[FFT.scala 34:12]
  assign _GEN_3847 = 7'h6 == cnt[6:0] ? $signed(32'shfd3b) : $signed(_GEN_3846); // @[FFT.scala 34:12]
  assign _GEN_3848 = 7'h7 == cnt[6:0] ? $signed(32'shfc3b) : $signed(_GEN_3847); // @[FFT.scala 34:12]
  assign _GEN_3849 = 7'h8 == cnt[6:0] ? $signed(32'shfb15) : $signed(_GEN_3848); // @[FFT.scala 34:12]
  assign _GEN_3850 = 7'h9 == cnt[6:0] ? $signed(32'shf9c8) : $signed(_GEN_3849); // @[FFT.scala 34:12]
  assign _GEN_3851 = 7'ha == cnt[6:0] ? $signed(32'shf854) : $signed(_GEN_3850); // @[FFT.scala 34:12]
  assign _GEN_3852 = 7'hb == cnt[6:0] ? $signed(32'shf6ba) : $signed(_GEN_3851); // @[FFT.scala 34:12]
  assign _GEN_3853 = 7'hc == cnt[6:0] ? $signed(32'shf4fa) : $signed(_GEN_3852); // @[FFT.scala 34:12]
  assign _GEN_3854 = 7'hd == cnt[6:0] ? $signed(32'shf314) : $signed(_GEN_3853); // @[FFT.scala 34:12]
  assign _GEN_3855 = 7'he == cnt[6:0] ? $signed(32'shf109) : $signed(_GEN_3854); // @[FFT.scala 34:12]
  assign _GEN_3856 = 7'hf == cnt[6:0] ? $signed(32'sheed9) : $signed(_GEN_3855); // @[FFT.scala 34:12]
  assign _GEN_3857 = 7'h10 == cnt[6:0] ? $signed(32'shec83) : $signed(_GEN_3856); // @[FFT.scala 34:12]
  assign _GEN_3858 = 7'h11 == cnt[6:0] ? $signed(32'shea0a) : $signed(_GEN_3857); // @[FFT.scala 34:12]
  assign _GEN_3859 = 7'h12 == cnt[6:0] ? $signed(32'she76c) : $signed(_GEN_3858); // @[FFT.scala 34:12]
  assign _GEN_3860 = 7'h13 == cnt[6:0] ? $signed(32'she4aa) : $signed(_GEN_3859); // @[FFT.scala 34:12]
  assign _GEN_3861 = 7'h14 == cnt[6:0] ? $signed(32'she1c6) : $signed(_GEN_3860); // @[FFT.scala 34:12]
  assign _GEN_3862 = 7'h15 == cnt[6:0] ? $signed(32'shdebe) : $signed(_GEN_3861); // @[FFT.scala 34:12]
  assign _GEN_3863 = 7'h16 == cnt[6:0] ? $signed(32'shdb94) : $signed(_GEN_3862); // @[FFT.scala 34:12]
  assign _GEN_3864 = 7'h17 == cnt[6:0] ? $signed(32'shd848) : $signed(_GEN_3863); // @[FFT.scala 34:12]
  assign _GEN_3865 = 7'h18 == cnt[6:0] ? $signed(32'shd4db) : $signed(_GEN_3864); // @[FFT.scala 34:12]
  assign _GEN_3866 = 7'h19 == cnt[6:0] ? $signed(32'shd14d) : $signed(_GEN_3865); // @[FFT.scala 34:12]
  assign _GEN_3867 = 7'h1a == cnt[6:0] ? $signed(32'shcd9f) : $signed(_GEN_3866); // @[FFT.scala 34:12]
  assign _GEN_3868 = 7'h1b == cnt[6:0] ? $signed(32'shc9d1) : $signed(_GEN_3867); // @[FFT.scala 34:12]
  assign _GEN_3869 = 7'h1c == cnt[6:0] ? $signed(32'shc5e4) : $signed(_GEN_3868); // @[FFT.scala 34:12]
  assign _GEN_3870 = 7'h1d == cnt[6:0] ? $signed(32'shc1d8) : $signed(_GEN_3869); // @[FFT.scala 34:12]
  assign _GEN_3871 = 7'h1e == cnt[6:0] ? $signed(32'shbdaf) : $signed(_GEN_3870); // @[FFT.scala 34:12]
  assign _GEN_3872 = 7'h1f == cnt[6:0] ? $signed(32'shb968) : $signed(_GEN_3871); // @[FFT.scala 34:12]
  assign _GEN_3873 = 7'h20 == cnt[6:0] ? $signed(32'shb505) : $signed(_GEN_3872); // @[FFT.scala 34:12]
  assign _GEN_3874 = 7'h21 == cnt[6:0] ? $signed(32'shb086) : $signed(_GEN_3873); // @[FFT.scala 34:12]
  assign _GEN_3875 = 7'h22 == cnt[6:0] ? $signed(32'shabeb) : $signed(_GEN_3874); // @[FFT.scala 34:12]
  assign _GEN_3876 = 7'h23 == cnt[6:0] ? $signed(32'sha736) : $signed(_GEN_3875); // @[FFT.scala 34:12]
  assign _GEN_3877 = 7'h24 == cnt[6:0] ? $signed(32'sha268) : $signed(_GEN_3876); // @[FFT.scala 34:12]
  assign _GEN_3878 = 7'h25 == cnt[6:0] ? $signed(32'sh9d80) : $signed(_GEN_3877); // @[FFT.scala 34:12]
  assign _GEN_3879 = 7'h26 == cnt[6:0] ? $signed(32'sh9880) : $signed(_GEN_3878); // @[FFT.scala 34:12]
  assign _GEN_3880 = 7'h27 == cnt[6:0] ? $signed(32'sh9368) : $signed(_GEN_3879); // @[FFT.scala 34:12]
  assign _GEN_3881 = 7'h28 == cnt[6:0] ? $signed(32'sh8e3a) : $signed(_GEN_3880); // @[FFT.scala 34:12]
  assign _GEN_3882 = 7'h29 == cnt[6:0] ? $signed(32'sh88f6) : $signed(_GEN_3881); // @[FFT.scala 34:12]
  assign _GEN_3883 = 7'h2a == cnt[6:0] ? $signed(32'sh839c) : $signed(_GEN_3882); // @[FFT.scala 34:12]
  assign _GEN_3884 = 7'h2b == cnt[6:0] ? $signed(32'sh7e2f) : $signed(_GEN_3883); // @[FFT.scala 34:12]
  assign _GEN_3885 = 7'h2c == cnt[6:0] ? $signed(32'sh78ad) : $signed(_GEN_3884); // @[FFT.scala 34:12]
  assign _GEN_3886 = 7'h2d == cnt[6:0] ? $signed(32'sh731a) : $signed(_GEN_3885); // @[FFT.scala 34:12]
  assign _GEN_3887 = 7'h2e == cnt[6:0] ? $signed(32'sh6d74) : $signed(_GEN_3886); // @[FFT.scala 34:12]
  assign _GEN_3888 = 7'h2f == cnt[6:0] ? $signed(32'sh67be) : $signed(_GEN_3887); // @[FFT.scala 34:12]
  assign _GEN_3889 = 7'h30 == cnt[6:0] ? $signed(32'sh61f8) : $signed(_GEN_3888); // @[FFT.scala 34:12]
  assign _GEN_3890 = 7'h31 == cnt[6:0] ? $signed(32'sh5c22) : $signed(_GEN_3889); // @[FFT.scala 34:12]
  assign _GEN_3891 = 7'h32 == cnt[6:0] ? $signed(32'sh563e) : $signed(_GEN_3890); // @[FFT.scala 34:12]
  assign _GEN_3892 = 7'h33 == cnt[6:0] ? $signed(32'sh504d) : $signed(_GEN_3891); // @[FFT.scala 34:12]
  assign _GEN_3893 = 7'h34 == cnt[6:0] ? $signed(32'sh4a50) : $signed(_GEN_3892); // @[FFT.scala 34:12]
  assign _GEN_3894 = 7'h35 == cnt[6:0] ? $signed(32'sh4447) : $signed(_GEN_3893); // @[FFT.scala 34:12]
  assign _GEN_3895 = 7'h36 == cnt[6:0] ? $signed(32'sh3e34) : $signed(_GEN_3894); // @[FFT.scala 34:12]
  assign _GEN_3896 = 7'h37 == cnt[6:0] ? $signed(32'sh3817) : $signed(_GEN_3895); // @[FFT.scala 34:12]
  assign _GEN_3897 = 7'h38 == cnt[6:0] ? $signed(32'sh31f1) : $signed(_GEN_3896); // @[FFT.scala 34:12]
  assign _GEN_3898 = 7'h39 == cnt[6:0] ? $signed(32'sh2bc4) : $signed(_GEN_3897); // @[FFT.scala 34:12]
  assign _GEN_3899 = 7'h3a == cnt[6:0] ? $signed(32'sh2590) : $signed(_GEN_3898); // @[FFT.scala 34:12]
  assign _GEN_3900 = 7'h3b == cnt[6:0] ? $signed(32'sh1f56) : $signed(_GEN_3899); // @[FFT.scala 34:12]
  assign _GEN_3901 = 7'h3c == cnt[6:0] ? $signed(32'sh1918) : $signed(_GEN_3900); // @[FFT.scala 34:12]
  assign _GEN_3902 = 7'h3d == cnt[6:0] ? $signed(32'sh12d5) : $signed(_GEN_3901); // @[FFT.scala 34:12]
  assign _GEN_3903 = 7'h3e == cnt[6:0] ? $signed(32'shc90) : $signed(_GEN_3902); // @[FFT.scala 34:12]
  assign _GEN_3904 = 7'h3f == cnt[6:0] ? $signed(32'sh648) : $signed(_GEN_3903); // @[FFT.scala 34:12]
  assign _GEN_3905 = 7'h40 == cnt[6:0] ? $signed(32'sh0) : $signed(_GEN_3904); // @[FFT.scala 34:12]
  assign _GEN_3906 = 7'h41 == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_3905); // @[FFT.scala 34:12]
  assign _GEN_3907 = 7'h42 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_3906); // @[FFT.scala 34:12]
  assign _GEN_3908 = 7'h43 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_3907); // @[FFT.scala 34:12]
  assign _GEN_3909 = 7'h44 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_3908); // @[FFT.scala 34:12]
  assign _GEN_3910 = 7'h45 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_3909); // @[FFT.scala 34:12]
  assign _GEN_3911 = 7'h46 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_3910); // @[FFT.scala 34:12]
  assign _GEN_3912 = 7'h47 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_3911); // @[FFT.scala 34:12]
  assign _GEN_3913 = 7'h48 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_3912); // @[FFT.scala 34:12]
  assign _GEN_3914 = 7'h49 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_3913); // @[FFT.scala 34:12]
  assign _GEN_3915 = 7'h4a == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_3914); // @[FFT.scala 34:12]
  assign _GEN_3916 = 7'h4b == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_3915); // @[FFT.scala 34:12]
  assign _GEN_3917 = 7'h4c == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_3916); // @[FFT.scala 34:12]
  assign _GEN_3918 = 7'h4d == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_3917); // @[FFT.scala 34:12]
  assign _GEN_3919 = 7'h4e == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_3918); // @[FFT.scala 34:12]
  assign _GEN_3920 = 7'h4f == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_3919); // @[FFT.scala 34:12]
  assign _GEN_3921 = 7'h50 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_3920); // @[FFT.scala 34:12]
  assign _GEN_3922 = 7'h51 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_3921); // @[FFT.scala 34:12]
  assign _GEN_3923 = 7'h52 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_3922); // @[FFT.scala 34:12]
  assign _GEN_3924 = 7'h53 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_3923); // @[FFT.scala 34:12]
  assign _GEN_3925 = 7'h54 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_3924); // @[FFT.scala 34:12]
  assign _GEN_3926 = 7'h55 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_3925); // @[FFT.scala 34:12]
  assign _GEN_3927 = 7'h56 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_3926); // @[FFT.scala 34:12]
  assign _GEN_3928 = 7'h57 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_3927); // @[FFT.scala 34:12]
  assign _GEN_3929 = 7'h58 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3928); // @[FFT.scala 34:12]
  assign _GEN_3930 = 7'h59 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_3929); // @[FFT.scala 34:12]
  assign _GEN_3931 = 7'h5a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_3930); // @[FFT.scala 34:12]
  assign _GEN_3932 = 7'h5b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_3931); // @[FFT.scala 34:12]
  assign _GEN_3933 = 7'h5c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_3932); // @[FFT.scala 34:12]
  assign _GEN_3934 = 7'h5d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_3933); // @[FFT.scala 34:12]
  assign _GEN_3935 = 7'h5e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_3934); // @[FFT.scala 34:12]
  assign _GEN_3936 = 7'h5f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_3935); // @[FFT.scala 34:12]
  assign _GEN_3937 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_3936); // @[FFT.scala 34:12]
  assign _GEN_3938 = 7'h61 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_3937); // @[FFT.scala 34:12]
  assign _GEN_3939 = 7'h62 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_3938); // @[FFT.scala 34:12]
  assign _GEN_3940 = 7'h63 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_3939); // @[FFT.scala 34:12]
  assign _GEN_3941 = 7'h64 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_3940); // @[FFT.scala 34:12]
  assign _GEN_3942 = 7'h65 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_3941); // @[FFT.scala 34:12]
  assign _GEN_3943 = 7'h66 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_3942); // @[FFT.scala 34:12]
  assign _GEN_3944 = 7'h67 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_3943); // @[FFT.scala 34:12]
  assign _GEN_3945 = 7'h68 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_3944); // @[FFT.scala 34:12]
  assign _GEN_3946 = 7'h69 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_3945); // @[FFT.scala 34:12]
  assign _GEN_3947 = 7'h6a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_3946); // @[FFT.scala 34:12]
  assign _GEN_3948 = 7'h6b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_3947); // @[FFT.scala 34:12]
  assign _GEN_3949 = 7'h6c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_3948); // @[FFT.scala 34:12]
  assign _GEN_3950 = 7'h6d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_3949); // @[FFT.scala 34:12]
  assign _GEN_3951 = 7'h6e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_3950); // @[FFT.scala 34:12]
  assign _GEN_3952 = 7'h6f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_3951); // @[FFT.scala 34:12]
  assign _GEN_3953 = 7'h70 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_3952); // @[FFT.scala 34:12]
  assign _GEN_3954 = 7'h71 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_3953); // @[FFT.scala 34:12]
  assign _GEN_3955 = 7'h72 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_3954); // @[FFT.scala 34:12]
  assign _GEN_3956 = 7'h73 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_3955); // @[FFT.scala 34:12]
  assign _GEN_3957 = 7'h74 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_3956); // @[FFT.scala 34:12]
  assign _GEN_3958 = 7'h75 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_3957); // @[FFT.scala 34:12]
  assign _GEN_3959 = 7'h76 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_3958); // @[FFT.scala 34:12]
  assign _GEN_3960 = 7'h77 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_3959); // @[FFT.scala 34:12]
  assign _GEN_3961 = 7'h78 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_3960); // @[FFT.scala 34:12]
  assign _GEN_3962 = 7'h79 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_3961); // @[FFT.scala 34:12]
  assign _GEN_3963 = 7'h7a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_3962); // @[FFT.scala 34:12]
  assign _GEN_3964 = 7'h7b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_3963); // @[FFT.scala 34:12]
  assign _GEN_3965 = 7'h7c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_3964); // @[FFT.scala 34:12]
  assign _GEN_3966 = 7'h7d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_3965); // @[FFT.scala 34:12]
  assign _GEN_3967 = 7'h7e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_3966); // @[FFT.scala 34:12]
  assign _GEN_3970 = 7'h1 == cnt[6:0] ? $signed(-32'sh648) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_3971 = 7'h2 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_3970); // @[FFT.scala 35:12]
  assign _GEN_3972 = 7'h3 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_3971); // @[FFT.scala 35:12]
  assign _GEN_3973 = 7'h4 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_3972); // @[FFT.scala 35:12]
  assign _GEN_3974 = 7'h5 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_3973); // @[FFT.scala 35:12]
  assign _GEN_3975 = 7'h6 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_3974); // @[FFT.scala 35:12]
  assign _GEN_3976 = 7'h7 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_3975); // @[FFT.scala 35:12]
  assign _GEN_3977 = 7'h8 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_3976); // @[FFT.scala 35:12]
  assign _GEN_3978 = 7'h9 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_3977); // @[FFT.scala 35:12]
  assign _GEN_3979 = 7'ha == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_3978); // @[FFT.scala 35:12]
  assign _GEN_3980 = 7'hb == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_3979); // @[FFT.scala 35:12]
  assign _GEN_3981 = 7'hc == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_3980); // @[FFT.scala 35:12]
  assign _GEN_3982 = 7'hd == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_3981); // @[FFT.scala 35:12]
  assign _GEN_3983 = 7'he == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_3982); // @[FFT.scala 35:12]
  assign _GEN_3984 = 7'hf == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_3983); // @[FFT.scala 35:12]
  assign _GEN_3985 = 7'h10 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_3984); // @[FFT.scala 35:12]
  assign _GEN_3986 = 7'h11 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_3985); // @[FFT.scala 35:12]
  assign _GEN_3987 = 7'h12 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_3986); // @[FFT.scala 35:12]
  assign _GEN_3988 = 7'h13 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_3987); // @[FFT.scala 35:12]
  assign _GEN_3989 = 7'h14 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_3988); // @[FFT.scala 35:12]
  assign _GEN_3990 = 7'h15 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_3989); // @[FFT.scala 35:12]
  assign _GEN_3991 = 7'h16 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_3990); // @[FFT.scala 35:12]
  assign _GEN_3992 = 7'h17 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_3991); // @[FFT.scala 35:12]
  assign _GEN_3993 = 7'h18 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3992); // @[FFT.scala 35:12]
  assign _GEN_3994 = 7'h19 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_3993); // @[FFT.scala 35:12]
  assign _GEN_3995 = 7'h1a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_3994); // @[FFT.scala 35:12]
  assign _GEN_3996 = 7'h1b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_3995); // @[FFT.scala 35:12]
  assign _GEN_3997 = 7'h1c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_3996); // @[FFT.scala 35:12]
  assign _GEN_3998 = 7'h1d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_3997); // @[FFT.scala 35:12]
  assign _GEN_3999 = 7'h1e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_3998); // @[FFT.scala 35:12]
  assign _GEN_4000 = 7'h1f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_3999); // @[FFT.scala 35:12]
  assign _GEN_4001 = 7'h20 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_4000); // @[FFT.scala 35:12]
  assign _GEN_4002 = 7'h21 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_4001); // @[FFT.scala 35:12]
  assign _GEN_4003 = 7'h22 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_4002); // @[FFT.scala 35:12]
  assign _GEN_4004 = 7'h23 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_4003); // @[FFT.scala 35:12]
  assign _GEN_4005 = 7'h24 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_4004); // @[FFT.scala 35:12]
  assign _GEN_4006 = 7'h25 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_4005); // @[FFT.scala 35:12]
  assign _GEN_4007 = 7'h26 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_4006); // @[FFT.scala 35:12]
  assign _GEN_4008 = 7'h27 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_4007); // @[FFT.scala 35:12]
  assign _GEN_4009 = 7'h28 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_4008); // @[FFT.scala 35:12]
  assign _GEN_4010 = 7'h29 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_4009); // @[FFT.scala 35:12]
  assign _GEN_4011 = 7'h2a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_4010); // @[FFT.scala 35:12]
  assign _GEN_4012 = 7'h2b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_4011); // @[FFT.scala 35:12]
  assign _GEN_4013 = 7'h2c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_4012); // @[FFT.scala 35:12]
  assign _GEN_4014 = 7'h2d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_4013); // @[FFT.scala 35:12]
  assign _GEN_4015 = 7'h2e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_4014); // @[FFT.scala 35:12]
  assign _GEN_4016 = 7'h2f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_4015); // @[FFT.scala 35:12]
  assign _GEN_4017 = 7'h30 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_4016); // @[FFT.scala 35:12]
  assign _GEN_4018 = 7'h31 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_4017); // @[FFT.scala 35:12]
  assign _GEN_4019 = 7'h32 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_4018); // @[FFT.scala 35:12]
  assign _GEN_4020 = 7'h33 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_4019); // @[FFT.scala 35:12]
  assign _GEN_4021 = 7'h34 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_4020); // @[FFT.scala 35:12]
  assign _GEN_4022 = 7'h35 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_4021); // @[FFT.scala 35:12]
  assign _GEN_4023 = 7'h36 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_4022); // @[FFT.scala 35:12]
  assign _GEN_4024 = 7'h37 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_4023); // @[FFT.scala 35:12]
  assign _GEN_4025 = 7'h38 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_4024); // @[FFT.scala 35:12]
  assign _GEN_4026 = 7'h39 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_4025); // @[FFT.scala 35:12]
  assign _GEN_4027 = 7'h3a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_4026); // @[FFT.scala 35:12]
  assign _GEN_4028 = 7'h3b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_4027); // @[FFT.scala 35:12]
  assign _GEN_4029 = 7'h3c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_4028); // @[FFT.scala 35:12]
  assign _GEN_4030 = 7'h3d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_4029); // @[FFT.scala 35:12]
  assign _GEN_4031 = 7'h3e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_4030); // @[FFT.scala 35:12]
  assign _GEN_4032 = 7'h3f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_4031); // @[FFT.scala 35:12]
  assign _GEN_4033 = 7'h40 == cnt[6:0] ? $signed(-32'sh10000) : $signed(_GEN_4032); // @[FFT.scala 35:12]
  assign _GEN_4034 = 7'h41 == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_4033); // @[FFT.scala 35:12]
  assign _GEN_4035 = 7'h42 == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_4034); // @[FFT.scala 35:12]
  assign _GEN_4036 = 7'h43 == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_4035); // @[FFT.scala 35:12]
  assign _GEN_4037 = 7'h44 == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_4036); // @[FFT.scala 35:12]
  assign _GEN_4038 = 7'h45 == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_4037); // @[FFT.scala 35:12]
  assign _GEN_4039 = 7'h46 == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_4038); // @[FFT.scala 35:12]
  assign _GEN_4040 = 7'h47 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_4039); // @[FFT.scala 35:12]
  assign _GEN_4041 = 7'h48 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_4040); // @[FFT.scala 35:12]
  assign _GEN_4042 = 7'h49 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_4041); // @[FFT.scala 35:12]
  assign _GEN_4043 = 7'h4a == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_4042); // @[FFT.scala 35:12]
  assign _GEN_4044 = 7'h4b == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_4043); // @[FFT.scala 35:12]
  assign _GEN_4045 = 7'h4c == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_4044); // @[FFT.scala 35:12]
  assign _GEN_4046 = 7'h4d == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_4045); // @[FFT.scala 35:12]
  assign _GEN_4047 = 7'h4e == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_4046); // @[FFT.scala 35:12]
  assign _GEN_4048 = 7'h4f == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_4047); // @[FFT.scala 35:12]
  assign _GEN_4049 = 7'h50 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_4048); // @[FFT.scala 35:12]
  assign _GEN_4050 = 7'h51 == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_4049); // @[FFT.scala 35:12]
  assign _GEN_4051 = 7'h52 == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_4050); // @[FFT.scala 35:12]
  assign _GEN_4052 = 7'h53 == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_4051); // @[FFT.scala 35:12]
  assign _GEN_4053 = 7'h54 == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_4052); // @[FFT.scala 35:12]
  assign _GEN_4054 = 7'h55 == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_4053); // @[FFT.scala 35:12]
  assign _GEN_4055 = 7'h56 == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_4054); // @[FFT.scala 35:12]
  assign _GEN_4056 = 7'h57 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_4055); // @[FFT.scala 35:12]
  assign _GEN_4057 = 7'h58 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_4056); // @[FFT.scala 35:12]
  assign _GEN_4058 = 7'h59 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_4057); // @[FFT.scala 35:12]
  assign _GEN_4059 = 7'h5a == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_4058); // @[FFT.scala 35:12]
  assign _GEN_4060 = 7'h5b == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_4059); // @[FFT.scala 35:12]
  assign _GEN_4061 = 7'h5c == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_4060); // @[FFT.scala 35:12]
  assign _GEN_4062 = 7'h5d == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_4061); // @[FFT.scala 35:12]
  assign _GEN_4063 = 7'h5e == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_4062); // @[FFT.scala 35:12]
  assign _GEN_4064 = 7'h5f == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_4063); // @[FFT.scala 35:12]
  assign _GEN_4065 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_4064); // @[FFT.scala 35:12]
  assign _GEN_4066 = 7'h61 == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_4065); // @[FFT.scala 35:12]
  assign _GEN_4067 = 7'h62 == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_4066); // @[FFT.scala 35:12]
  assign _GEN_4068 = 7'h63 == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_4067); // @[FFT.scala 35:12]
  assign _GEN_4069 = 7'h64 == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_4068); // @[FFT.scala 35:12]
  assign _GEN_4070 = 7'h65 == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_4069); // @[FFT.scala 35:12]
  assign _GEN_4071 = 7'h66 == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_4070); // @[FFT.scala 35:12]
  assign _GEN_4072 = 7'h67 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_4071); // @[FFT.scala 35:12]
  assign _GEN_4073 = 7'h68 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4072); // @[FFT.scala 35:12]
  assign _GEN_4074 = 7'h69 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_4073); // @[FFT.scala 35:12]
  assign _GEN_4075 = 7'h6a == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_4074); // @[FFT.scala 35:12]
  assign _GEN_4076 = 7'h6b == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_4075); // @[FFT.scala 35:12]
  assign _GEN_4077 = 7'h6c == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_4076); // @[FFT.scala 35:12]
  assign _GEN_4078 = 7'h6d == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_4077); // @[FFT.scala 35:12]
  assign _GEN_4079 = 7'h6e == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_4078); // @[FFT.scala 35:12]
  assign _GEN_4080 = 7'h6f == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_4079); // @[FFT.scala 35:12]
  assign _GEN_4081 = 7'h70 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_4080); // @[FFT.scala 35:12]
  assign _GEN_4082 = 7'h71 == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_4081); // @[FFT.scala 35:12]
  assign _GEN_4083 = 7'h72 == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_4082); // @[FFT.scala 35:12]
  assign _GEN_4084 = 7'h73 == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_4083); // @[FFT.scala 35:12]
  assign _GEN_4085 = 7'h74 == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_4084); // @[FFT.scala 35:12]
  assign _GEN_4086 = 7'h75 == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_4085); // @[FFT.scala 35:12]
  assign _GEN_4087 = 7'h76 == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_4086); // @[FFT.scala 35:12]
  assign _GEN_4088 = 7'h77 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_4087); // @[FFT.scala 35:12]
  assign _GEN_4089 = 7'h78 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_4088); // @[FFT.scala 35:12]
  assign _GEN_4090 = 7'h79 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_4089); // @[FFT.scala 35:12]
  assign _GEN_4091 = 7'h7a == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_4090); // @[FFT.scala 35:12]
  assign _GEN_4092 = 7'h7b == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_4091); // @[FFT.scala 35:12]
  assign _GEN_4093 = 7'h7c == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_4092); // @[FFT.scala 35:12]
  assign _GEN_4094 = 7'h7d == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_4093); // @[FFT.scala 35:12]
  assign _GEN_4095 = 7'h7e == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_4094); // @[FFT.scala 35:12]
  assign _GEN_4482 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_4483 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_4482); // @[FFT.scala 34:12]
  assign _GEN_4484 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_4483); // @[FFT.scala 34:12]
  assign _GEN_4485 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_4484); // @[FFT.scala 34:12]
  assign _GEN_4486 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_4485); // @[FFT.scala 34:12]
  assign _GEN_4487 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_4486); // @[FFT.scala 34:12]
  assign _GEN_4488 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_4487); // @[FFT.scala 34:12]
  assign _GEN_4489 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_4488); // @[FFT.scala 34:12]
  assign _GEN_4490 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_4489); // @[FFT.scala 34:12]
  assign _GEN_4491 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_4490); // @[FFT.scala 34:12]
  assign _GEN_4492 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_4491); // @[FFT.scala 34:12]
  assign _GEN_4493 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_4492); // @[FFT.scala 34:12]
  assign _GEN_4494 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_4493); // @[FFT.scala 34:12]
  assign _GEN_4495 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_4494); // @[FFT.scala 34:12]
  assign _GEN_4496 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_4495); // @[FFT.scala 34:12]
  assign _GEN_4497 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_4496); // @[FFT.scala 34:12]
  assign _GEN_4498 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_4497); // @[FFT.scala 34:12]
  assign _GEN_4499 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_4498); // @[FFT.scala 34:12]
  assign _GEN_4500 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_4499); // @[FFT.scala 34:12]
  assign _GEN_4501 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_4500); // @[FFT.scala 34:12]
  assign _GEN_4502 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_4501); // @[FFT.scala 34:12]
  assign _GEN_4503 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_4502); // @[FFT.scala 34:12]
  assign _GEN_4504 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_4503); // @[FFT.scala 34:12]
  assign _GEN_4505 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_4504); // @[FFT.scala 34:12]
  assign _GEN_4506 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_4505); // @[FFT.scala 34:12]
  assign _GEN_4507 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_4506); // @[FFT.scala 34:12]
  assign _GEN_4508 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_4507); // @[FFT.scala 34:12]
  assign _GEN_4509 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_4508); // @[FFT.scala 34:12]
  assign _GEN_4510 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_4509); // @[FFT.scala 34:12]
  assign _GEN_4511 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_4510); // @[FFT.scala 34:12]
  assign _GEN_4512 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_4511); // @[FFT.scala 34:12]
  assign _GEN_4513 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_4512); // @[FFT.scala 34:12]
  assign _GEN_4514 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_4513); // @[FFT.scala 34:12]
  assign _GEN_4515 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_4514); // @[FFT.scala 34:12]
  assign _GEN_4516 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_4515); // @[FFT.scala 34:12]
  assign _GEN_4517 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_4516); // @[FFT.scala 34:12]
  assign _GEN_4518 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_4517); // @[FFT.scala 34:12]
  assign _GEN_4519 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_4518); // @[FFT.scala 34:12]
  assign _GEN_4520 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_4519); // @[FFT.scala 34:12]
  assign _GEN_4521 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_4520); // @[FFT.scala 34:12]
  assign _GEN_4522 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_4521); // @[FFT.scala 34:12]
  assign _GEN_4523 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_4522); // @[FFT.scala 34:12]
  assign _GEN_4524 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_4523); // @[FFT.scala 34:12]
  assign _GEN_4525 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4524); // @[FFT.scala 34:12]
  assign _GEN_4526 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_4525); // @[FFT.scala 34:12]
  assign _GEN_4527 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_4526); // @[FFT.scala 34:12]
  assign _GEN_4528 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_4527); // @[FFT.scala 34:12]
  assign _GEN_4529 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_4528); // @[FFT.scala 34:12]
  assign _GEN_4530 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_4529); // @[FFT.scala 34:12]
  assign _GEN_4531 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_4530); // @[FFT.scala 34:12]
  assign _GEN_4532 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_4531); // @[FFT.scala 34:12]
  assign _GEN_4533 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_4532); // @[FFT.scala 34:12]
  assign _GEN_4534 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_4533); // @[FFT.scala 34:12]
  assign _GEN_4535 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_4534); // @[FFT.scala 34:12]
  assign _GEN_4536 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_4535); // @[FFT.scala 34:12]
  assign _GEN_4537 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_4536); // @[FFT.scala 34:12]
  assign _GEN_4538 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_4537); // @[FFT.scala 34:12]
  assign _GEN_4539 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_4538); // @[FFT.scala 34:12]
  assign _GEN_4540 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_4539); // @[FFT.scala 34:12]
  assign _GEN_4541 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_4540); // @[FFT.scala 34:12]
  assign _GEN_4542 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_4541); // @[FFT.scala 34:12]
  assign _GEN_4543 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_4542); // @[FFT.scala 34:12]
  assign _GEN_4546 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_4547 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_4546); // @[FFT.scala 35:12]
  assign _GEN_4548 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_4547); // @[FFT.scala 35:12]
  assign _GEN_4549 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_4548); // @[FFT.scala 35:12]
  assign _GEN_4550 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_4549); // @[FFT.scala 35:12]
  assign _GEN_4551 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_4550); // @[FFT.scala 35:12]
  assign _GEN_4552 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_4551); // @[FFT.scala 35:12]
  assign _GEN_4553 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_4552); // @[FFT.scala 35:12]
  assign _GEN_4554 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_4553); // @[FFT.scala 35:12]
  assign _GEN_4555 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_4554); // @[FFT.scala 35:12]
  assign _GEN_4556 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_4555); // @[FFT.scala 35:12]
  assign _GEN_4557 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4556); // @[FFT.scala 35:12]
  assign _GEN_4558 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_4557); // @[FFT.scala 35:12]
  assign _GEN_4559 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_4558); // @[FFT.scala 35:12]
  assign _GEN_4560 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_4559); // @[FFT.scala 35:12]
  assign _GEN_4561 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_4560); // @[FFT.scala 35:12]
  assign _GEN_4562 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_4561); // @[FFT.scala 35:12]
  assign _GEN_4563 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_4562); // @[FFT.scala 35:12]
  assign _GEN_4564 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_4563); // @[FFT.scala 35:12]
  assign _GEN_4565 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_4564); // @[FFT.scala 35:12]
  assign _GEN_4566 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_4565); // @[FFT.scala 35:12]
  assign _GEN_4567 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_4566); // @[FFT.scala 35:12]
  assign _GEN_4568 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_4567); // @[FFT.scala 35:12]
  assign _GEN_4569 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_4568); // @[FFT.scala 35:12]
  assign _GEN_4570 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_4569); // @[FFT.scala 35:12]
  assign _GEN_4571 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_4570); // @[FFT.scala 35:12]
  assign _GEN_4572 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_4571); // @[FFT.scala 35:12]
  assign _GEN_4573 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_4572); // @[FFT.scala 35:12]
  assign _GEN_4574 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_4573); // @[FFT.scala 35:12]
  assign _GEN_4575 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_4574); // @[FFT.scala 35:12]
  assign _GEN_4576 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_4575); // @[FFT.scala 35:12]
  assign _GEN_4577 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_4576); // @[FFT.scala 35:12]
  assign _GEN_4578 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_4577); // @[FFT.scala 35:12]
  assign _GEN_4579 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_4578); // @[FFT.scala 35:12]
  assign _GEN_4580 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_4579); // @[FFT.scala 35:12]
  assign _GEN_4581 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_4580); // @[FFT.scala 35:12]
  assign _GEN_4582 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_4581); // @[FFT.scala 35:12]
  assign _GEN_4583 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_4582); // @[FFT.scala 35:12]
  assign _GEN_4584 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_4583); // @[FFT.scala 35:12]
  assign _GEN_4585 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_4584); // @[FFT.scala 35:12]
  assign _GEN_4586 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_4585); // @[FFT.scala 35:12]
  assign _GEN_4587 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_4586); // @[FFT.scala 35:12]
  assign _GEN_4588 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_4587); // @[FFT.scala 35:12]
  assign _GEN_4589 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_4588); // @[FFT.scala 35:12]
  assign _GEN_4590 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_4589); // @[FFT.scala 35:12]
  assign _GEN_4591 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_4590); // @[FFT.scala 35:12]
  assign _GEN_4592 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_4591); // @[FFT.scala 35:12]
  assign _GEN_4593 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_4592); // @[FFT.scala 35:12]
  assign _GEN_4594 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_4593); // @[FFT.scala 35:12]
  assign _GEN_4595 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_4594); // @[FFT.scala 35:12]
  assign _GEN_4596 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_4595); // @[FFT.scala 35:12]
  assign _GEN_4597 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4596); // @[FFT.scala 35:12]
  assign _GEN_4598 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_4597); // @[FFT.scala 35:12]
  assign _GEN_4599 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_4598); // @[FFT.scala 35:12]
  assign _GEN_4600 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_4599); // @[FFT.scala 35:12]
  assign _GEN_4601 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_4600); // @[FFT.scala 35:12]
  assign _GEN_4602 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_4601); // @[FFT.scala 35:12]
  assign _GEN_4603 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_4602); // @[FFT.scala 35:12]
  assign _GEN_4604 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_4603); // @[FFT.scala 35:12]
  assign _GEN_4605 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_4604); // @[FFT.scala 35:12]
  assign _GEN_4606 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_4605); // @[FFT.scala 35:12]
  assign _GEN_4607 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_4606); // @[FFT.scala 35:12]
  assign _GEN_4802 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_4803 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_4802); // @[FFT.scala 34:12]
  assign _GEN_4804 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_4803); // @[FFT.scala 34:12]
  assign _GEN_4805 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_4804); // @[FFT.scala 34:12]
  assign _GEN_4806 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_4805); // @[FFT.scala 34:12]
  assign _GEN_4807 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_4806); // @[FFT.scala 34:12]
  assign _GEN_4808 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_4807); // @[FFT.scala 34:12]
  assign _GEN_4809 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_4808); // @[FFT.scala 34:12]
  assign _GEN_4810 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_4809); // @[FFT.scala 34:12]
  assign _GEN_4811 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_4810); // @[FFT.scala 34:12]
  assign _GEN_4812 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_4811); // @[FFT.scala 34:12]
  assign _GEN_4813 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_4812); // @[FFT.scala 34:12]
  assign _GEN_4814 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_4813); // @[FFT.scala 34:12]
  assign _GEN_4815 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_4814); // @[FFT.scala 34:12]
  assign _GEN_4816 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_4815); // @[FFT.scala 34:12]
  assign _GEN_4817 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_4816); // @[FFT.scala 34:12]
  assign _GEN_4818 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_4817); // @[FFT.scala 34:12]
  assign _GEN_4819 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_4818); // @[FFT.scala 34:12]
  assign _GEN_4820 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_4819); // @[FFT.scala 34:12]
  assign _GEN_4821 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_4820); // @[FFT.scala 34:12]
  assign _GEN_4822 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_4821); // @[FFT.scala 34:12]
  assign _GEN_4823 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4822); // @[FFT.scala 34:12]
  assign _GEN_4824 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_4823); // @[FFT.scala 34:12]
  assign _GEN_4825 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_4824); // @[FFT.scala 34:12]
  assign _GEN_4826 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_4825); // @[FFT.scala 34:12]
  assign _GEN_4827 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_4826); // @[FFT.scala 34:12]
  assign _GEN_4828 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_4827); // @[FFT.scala 34:12]
  assign _GEN_4829 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_4828); // @[FFT.scala 34:12]
  assign _GEN_4830 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_4829); // @[FFT.scala 34:12]
  assign _GEN_4831 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_4830); // @[FFT.scala 34:12]
  assign _GEN_4834 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_4835 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_4834); // @[FFT.scala 35:12]
  assign _GEN_4836 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_4835); // @[FFT.scala 35:12]
  assign _GEN_4837 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_4836); // @[FFT.scala 35:12]
  assign _GEN_4838 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_4837); // @[FFT.scala 35:12]
  assign _GEN_4839 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4838); // @[FFT.scala 35:12]
  assign _GEN_4840 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_4839); // @[FFT.scala 35:12]
  assign _GEN_4841 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_4840); // @[FFT.scala 35:12]
  assign _GEN_4842 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_4841); // @[FFT.scala 35:12]
  assign _GEN_4843 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_4842); // @[FFT.scala 35:12]
  assign _GEN_4844 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_4843); // @[FFT.scala 35:12]
  assign _GEN_4845 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_4844); // @[FFT.scala 35:12]
  assign _GEN_4846 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_4845); // @[FFT.scala 35:12]
  assign _GEN_4847 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_4846); // @[FFT.scala 35:12]
  assign _GEN_4848 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_4847); // @[FFT.scala 35:12]
  assign _GEN_4849 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_4848); // @[FFT.scala 35:12]
  assign _GEN_4850 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_4849); // @[FFT.scala 35:12]
  assign _GEN_4851 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_4850); // @[FFT.scala 35:12]
  assign _GEN_4852 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_4851); // @[FFT.scala 35:12]
  assign _GEN_4853 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_4852); // @[FFT.scala 35:12]
  assign _GEN_4854 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_4853); // @[FFT.scala 35:12]
  assign _GEN_4855 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_4854); // @[FFT.scala 35:12]
  assign _GEN_4856 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_4855); // @[FFT.scala 35:12]
  assign _GEN_4857 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_4856); // @[FFT.scala 35:12]
  assign _GEN_4858 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_4857); // @[FFT.scala 35:12]
  assign _GEN_4859 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4858); // @[FFT.scala 35:12]
  assign _GEN_4860 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_4859); // @[FFT.scala 35:12]
  assign _GEN_4861 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_4860); // @[FFT.scala 35:12]
  assign _GEN_4862 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_4861); // @[FFT.scala 35:12]
  assign _GEN_4863 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_4862); // @[FFT.scala 35:12]
  assign _GEN_4962 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_4963 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_4962); // @[FFT.scala 34:12]
  assign _GEN_4964 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_4963); // @[FFT.scala 34:12]
  assign _GEN_4965 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_4964); // @[FFT.scala 34:12]
  assign _GEN_4966 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_4965); // @[FFT.scala 34:12]
  assign _GEN_4967 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_4966); // @[FFT.scala 34:12]
  assign _GEN_4968 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_4967); // @[FFT.scala 34:12]
  assign _GEN_4969 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_4968); // @[FFT.scala 34:12]
  assign _GEN_4970 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_4969); // @[FFT.scala 34:12]
  assign _GEN_4971 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_4970); // @[FFT.scala 34:12]
  assign _GEN_4972 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4971); // @[FFT.scala 34:12]
  assign _GEN_4973 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_4972); // @[FFT.scala 34:12]
  assign _GEN_4974 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_4973); // @[FFT.scala 34:12]
  assign _GEN_4975 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_4974); // @[FFT.scala 34:12]
  assign _GEN_4978 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_4979 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_4978); // @[FFT.scala 35:12]
  assign _GEN_4980 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4979); // @[FFT.scala 35:12]
  assign _GEN_4981 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_4980); // @[FFT.scala 35:12]
  assign _GEN_4982 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_4981); // @[FFT.scala 35:12]
  assign _GEN_4983 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_4982); // @[FFT.scala 35:12]
  assign _GEN_4984 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_4983); // @[FFT.scala 35:12]
  assign _GEN_4985 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_4984); // @[FFT.scala 35:12]
  assign _GEN_4986 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_4985); // @[FFT.scala 35:12]
  assign _GEN_4987 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_4986); // @[FFT.scala 35:12]
  assign _GEN_4988 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_4987); // @[FFT.scala 35:12]
  assign _GEN_4989 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_4988); // @[FFT.scala 35:12]
  assign _GEN_4990 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_4989); // @[FFT.scala 35:12]
  assign _GEN_4991 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_4990); // @[FFT.scala 35:12]
  assign _GEN_5042 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_5043 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_5042); // @[FFT.scala 34:12]
  assign _GEN_5044 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_5043); // @[FFT.scala 34:12]
  assign _GEN_5045 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_5044); // @[FFT.scala 34:12]
  assign _GEN_5046 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_5045); // @[FFT.scala 34:12]
  assign _GEN_5047 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_5046); // @[FFT.scala 34:12]
  assign _GEN_5050 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_5051 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_5050); // @[FFT.scala 35:12]
  assign _GEN_5052 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_5051); // @[FFT.scala 35:12]
  assign _GEN_5053 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_5052); // @[FFT.scala 35:12]
  assign _GEN_5054 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_5053); // @[FFT.scala 35:12]
  assign _GEN_5055 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_5054); // @[FFT.scala 35:12]
  assign _GEN_5082 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_5083 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_5082); // @[FFT.scala 34:12]
  assign _GEN_5086 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_5087 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_5086); // @[FFT.scala 35:12]
  assign io_dOut1_re = _T_1752_re; // @[FFT.scala 85:12]
  assign io_dOut1_im = _T_1752_im; // @[FFT.scala 85:12]
  assign io_dOut2_re = _T_1753_re; // @[FFT.scala 86:12]
  assign io_dOut2_im = _T_1753_im; // @[FFT.scala 86:12]
  assign io_dout_valid = cntD1 == 10'h3ff; // @[FFT.scala 91:19]
  assign Butterfly_io_in1_re = _T_672_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_672_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = io_dIn_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = 9'h1ff == cnt[8:0] ? $signed(-32'shffff) : $signed(_GEN_511); // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = 9'h1ff == cnt[8:0] ? $signed(-32'sh192) : $signed(_GEN_1023); // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_930_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_930_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cnt[8]; // @[Butterfly.scala 113:17]
  assign Butterfly_1_io_in1_re = _T_1191_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_1191_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = 8'hff == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_2815); // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = 8'hff == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_3071); // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_1321_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_1321_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cnt[7]; // @[Butterfly.scala 113:17]
  assign Butterfly_2_io_in1_re = _T_1454_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_1454_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = 7'h7f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_3967); // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = 7'h7f == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_4095); // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_1520_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_1520_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cnt[6]; // @[Butterfly.scala 113:17]
  assign Butterfly_3_io_in1_re = _T_1589_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_1589_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_4543); // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_4607); // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_1623_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_1623_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cnt[5]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_1660_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_1660_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_4831); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_4863); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_1678_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_1678_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cnt[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_1699_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_1699_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_4975); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_4991); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_1709_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_1709_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cnt[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_1722_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_1722_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_5047); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_5055); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_1728_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_1728_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cnt[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_7_io_in1_re = _T_1737_re; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in1_im = _T_1737_im; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_5083); // @[Butterfly.scala 92:16]
  assign Butterfly_7_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_5087); // @[Butterfly.scala 92:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in2_re = _T_1741_re; // @[Butterfly.scala 112:17]
  assign Switch_7_io_in2_im = _T_1741_im; // @[Butterfly.scala 112:17]
  assign Switch_7_io_sel = cnt[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_8_io_in1_re = _T_1748_re; // @[Butterfly.scala 90:17]
  assign Butterfly_8_io_in1_im = _T_1748_im; // @[Butterfly.scala 90:17]
  assign Butterfly_8_io_in2_re = Switch_7_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_8_io_in2_im = Switch_7_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_8_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_8_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_8_io_in1_re = Butterfly_8_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_8_io_in1_im = Butterfly_8_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_8_io_in2_re = _T_1751_re; // @[Butterfly.scala 112:17]
  assign Switch_8_io_in2_im = _T_1751_im; // @[Butterfly.scala 112:17]
  assign Switch_8_io_sel = cnt[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_8_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_8_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_8_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_8_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntD1 = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_161_re = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_161_im = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_162_re = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_162_im = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_163_re = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_163_im = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_164_re = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_164_im = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_165_re = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_165_im = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_166_re = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_166_im = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_167_re = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_167_im = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_168_re = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_168_im = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_169_re = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_169_im = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_170_re = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_170_im = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_171_re = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_171_im = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_172_re = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_172_im = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_173_re = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_173_im = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_174_re = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_174_im = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_175_re = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_175_im = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_176_re = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_176_im = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_177_re = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_177_im = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_178_re = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_178_im = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_179_re = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_179_im = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_180_re = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_180_im = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_181_re = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_181_im = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_182_re = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_182_im = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_183_re = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_183_im = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_184_re = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_184_im = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_185_re = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_185_im = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_186_re = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_186_im = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_187_re = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_187_im = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_188_re = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_188_im = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_189_re = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_189_im = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_190_re = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_190_im = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_191_re = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_191_im = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_192_re = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_192_im = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_193_re = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_193_im = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_194_re = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_194_im = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_195_re = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_195_im = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_196_re = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_196_im = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_197_re = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_197_im = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_198_re = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_198_im = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_199_re = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_199_im = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_200_re = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_200_im = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_201_re = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_201_im = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_202_re = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_202_im = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_203_re = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_203_im = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_204_re = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_204_im = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_205_re = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_205_im = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_206_re = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_206_im = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_207_re = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_207_im = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_208_re = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_208_im = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_209_re = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_209_im = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_210_re = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_210_im = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_211_re = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_211_im = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_212_re = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_212_im = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_213_re = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_213_im = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_214_re = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_214_im = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_215_re = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_215_im = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_216_re = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_216_im = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_217_re = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_217_im = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_218_re = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_218_im = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_219_re = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_219_im = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_220_re = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_220_im = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_221_re = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_221_im = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_222_re = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_222_im = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_223_re = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_223_im = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_224_re = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_224_im = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_225_re = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_225_im = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_226_re = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_226_im = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_227_re = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_227_im = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_228_re = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_228_im = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_229_re = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_229_im = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_230_re = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_230_im = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_231_re = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_231_im = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_232_re = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_232_im = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_233_re = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_233_im = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_234_re = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_234_im = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_235_re = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_235_im = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_236_re = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_236_im = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_237_re = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_237_im = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_238_re = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_238_im = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_239_re = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_239_im = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_240_re = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_240_im = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_241_re = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_241_im = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_242_re = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_242_im = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_243_re = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_243_im = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_244_re = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_244_im = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_245_re = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_245_im = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_246_re = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_246_im = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_247_re = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_247_im = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_248_re = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_248_im = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_249_re = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_249_im = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_250_re = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_250_im = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_251_re = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_251_im = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_252_re = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_252_im = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_253_re = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_253_im = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_254_re = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_254_im = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_255_re = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_255_im = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_256_re = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_256_im = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_257_re = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_257_im = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_258_re = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_258_im = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_259_re = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_259_im = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_260_re = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_260_im = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_261_re = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_261_im = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_262_re = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_262_im = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_263_re = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_263_im = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_264_re = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_264_im = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_265_re = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_265_im = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_266_re = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_266_im = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_267_re = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_267_im = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_268_re = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_268_im = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_269_re = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_269_im = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_270_re = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_270_im = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_271_re = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_271_im = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_272_re = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_272_im = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_273_re = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_273_im = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_274_re = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_274_im = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_275_re = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_275_im = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_276_re = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_276_im = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_277_re = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_277_im = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_278_re = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_278_im = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_279_re = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_279_im = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_280_re = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_280_im = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_281_re = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_281_im = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_282_re = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_282_im = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_283_re = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_283_im = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_284_re = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_284_im = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_285_re = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_285_im = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_286_re = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_286_im = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_287_re = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_287_im = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_288_re = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_288_im = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_289_re = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_289_im = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_290_re = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_290_im = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_291_re = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_291_im = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_292_re = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_292_im = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_293_re = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_293_im = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_294_re = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_294_im = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_295_re = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_295_im = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_296_re = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_296_im = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_297_re = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_297_im = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_298_re = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_298_im = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_299_re = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_299_im = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_300_re = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_300_im = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_301_re = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_301_im = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_302_re = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_302_im = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_303_re = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_303_im = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_304_re = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_304_im = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_305_re = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_305_im = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_306_re = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_306_im = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_307_re = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_307_im = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_308_re = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_308_im = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_309_re = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_309_im = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_310_re = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_310_im = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_311_re = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_311_im = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_312_re = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_312_im = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_313_re = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_313_im = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_314_re = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_314_im = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_315_re = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_315_im = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_316_re = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_316_im = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_317_re = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_317_im = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_318_re = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_318_im = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_319_re = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_319_im = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_320_re = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_320_im = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_321_re = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_321_im = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_322_re = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_322_im = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_323_re = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_323_im = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_324_re = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_324_im = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_325_re = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_325_im = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_326_re = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_326_im = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_327_re = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_327_im = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_328_re = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_328_im = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_329_re = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_329_im = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_330_re = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_330_im = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_331_re = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_331_im = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_332_re = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_332_im = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_333_re = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_333_im = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_334_re = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_334_im = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_335_re = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_335_im = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_336_re = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_336_im = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_337_re = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_337_im = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_338_re = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_338_im = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_339_re = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_339_im = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_340_re = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_340_im = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_341_re = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_341_im = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_342_re = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_342_im = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_343_re = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_343_im = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_344_re = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_344_im = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_345_re = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_345_im = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_346_re = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_346_im = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_347_re = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_347_im = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_348_re = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_348_im = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_349_re = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_349_im = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_350_re = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_350_im = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_351_re = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_351_im = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_352_re = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_352_im = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_353_re = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_353_im = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_354_re = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_354_im = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_355_re = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_355_im = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_356_re = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_356_im = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_357_re = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_357_im = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_358_re = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_358_im = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_359_re = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_359_im = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_360_re = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_360_im = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_361_re = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_361_im = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_362_re = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_362_im = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_363_re = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_363_im = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_364_re = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_364_im = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_365_re = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_365_im = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_366_re = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_366_im = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_367_re = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_367_im = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_368_re = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_368_im = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_369_re = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_369_im = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_370_re = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_370_im = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_371_re = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_371_im = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_372_re = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_372_im = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_373_re = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_373_im = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_374_re = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_374_im = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_375_re = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_375_im = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_376_re = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_376_im = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_377_re = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_377_im = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_378_re = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_378_im = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_379_re = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_379_im = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_380_re = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_380_im = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_381_re = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_381_im = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_382_re = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_382_im = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_383_re = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_383_im = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_384_re = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_384_im = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_385_re = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_385_im = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_386_re = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_386_im = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_387_re = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_387_im = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_388_re = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_388_im = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_389_re = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_389_im = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_390_re = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_390_im = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_391_re = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_391_im = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_392_re = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_392_im = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_393_re = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_393_im = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_394_re = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_394_im = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_395_re = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_395_im = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_396_re = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_396_im = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_397_re = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_397_im = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_398_re = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_398_im = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_399_re = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_399_im = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_400_re = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_400_im = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_401_re = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_401_im = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_402_re = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_402_im = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_403_re = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_403_im = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_404_re = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_404_im = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_405_re = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_405_im = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_406_re = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_406_im = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_407_re = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_407_im = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_408_re = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_408_im = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_409_re = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_409_im = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_410_re = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_410_im = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_411_re = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_411_im = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_412_re = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_412_im = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_413_re = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_413_im = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_414_re = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_414_im = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_415_re = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_415_im = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_416_re = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_416_im = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_417_re = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_417_im = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_418_re = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_418_im = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_419_re = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_419_im = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_420_re = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_420_im = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_421_re = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_421_im = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_422_re = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_422_im = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_423_re = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_423_im = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_424_re = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_424_im = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_425_re = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_425_im = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_426_re = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_426_im = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_427_re = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_427_im = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_428_re = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_428_im = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_429_re = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_429_im = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_430_re = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_430_im = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_431_re = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_431_im = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_432_re = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_432_im = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_433_re = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_433_im = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_434_re = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_434_im = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_435_re = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_435_im = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_436_re = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_436_im = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_437_re = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_437_im = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_438_re = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_438_im = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_439_re = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_439_im = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_440_re = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_440_im = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_441_re = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_441_im = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_442_re = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_442_im = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_443_re = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_443_im = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_444_re = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_444_im = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_445_re = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_445_im = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_446_re = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_446_im = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_447_re = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_447_im = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_448_re = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_448_im = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_449_re = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_449_im = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_450_re = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_450_im = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_451_re = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_451_im = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_452_re = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_452_im = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_453_re = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_453_im = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_454_re = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_454_im = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_455_re = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_455_im = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_456_re = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_456_im = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_457_re = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_457_im = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_458_re = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_458_im = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_459_re = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_459_im = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_460_re = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_460_im = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_461_re = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_461_im = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_462_re = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_462_im = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_463_re = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_463_im = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_464_re = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_464_im = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_465_re = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_465_im = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_466_re = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_466_im = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_467_re = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_467_im = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_468_re = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_468_im = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_469_re = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_469_im = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_470_re = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_470_im = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_471_re = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_471_im = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_472_re = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_472_im = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_473_re = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_473_im = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_474_re = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_474_im = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_475_re = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_475_im = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_476_re = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_476_im = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_477_re = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_477_im = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_478_re = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_478_im = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_479_re = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_479_im = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_480_re = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_480_im = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_481_re = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_481_im = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_482_re = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_482_im = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_483_re = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_483_im = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_484_re = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_484_im = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_485_re = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_485_im = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_486_re = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_486_im = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_487_re = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_487_im = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_488_re = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_488_im = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_489_re = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_489_im = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_490_re = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_490_im = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_491_re = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_491_im = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_492_re = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_492_im = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_493_re = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_493_im = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_494_re = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_494_im = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_495_re = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_495_im = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_496_re = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_496_im = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_497_re = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_497_im = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_498_re = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_498_im = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_499_re = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_499_im = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_500_re = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_500_im = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_501_re = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_501_im = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_502_re = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_502_im = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_503_re = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_503_im = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_504_re = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_504_im = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_505_re = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_505_im = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_506_re = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_506_im = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_507_re = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_507_im = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_508_re = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_508_im = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_509_re = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_509_im = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_510_re = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_510_im = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_511_re = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_511_im = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_512_re = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_512_im = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_513_re = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_513_im = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_514_re = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_514_im = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_515_re = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_515_im = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_516_re = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_516_im = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_517_re = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_517_im = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_518_re = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_518_im = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_519_re = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_519_im = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_520_re = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_520_im = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_521_re = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_521_im = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_522_re = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_522_im = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_523_re = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_523_im = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_524_re = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_524_im = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_525_re = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_525_im = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_526_re = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_526_im = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_527_re = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_527_im = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_528_re = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_528_im = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_529_re = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_529_im = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_530_re = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_530_im = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_531_re = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_531_im = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_532_re = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_532_im = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_533_re = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_533_im = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_534_re = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_534_im = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_535_re = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_535_im = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_536_re = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_536_im = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_537_re = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_537_im = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_538_re = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_538_im = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_539_re = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_539_im = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_540_re = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_540_im = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_541_re = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_541_im = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_542_re = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_542_im = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_543_re = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_543_im = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_544_re = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_544_im = _RAND_769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_545_re = _RAND_770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_545_im = _RAND_771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_546_re = _RAND_772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_546_im = _RAND_773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_547_re = _RAND_774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_547_im = _RAND_775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_548_re = _RAND_776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_548_im = _RAND_777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_549_re = _RAND_778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_549_im = _RAND_779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_550_re = _RAND_780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_550_im = _RAND_781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_551_re = _RAND_782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_551_im = _RAND_783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_552_re = _RAND_784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_552_im = _RAND_785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_553_re = _RAND_786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_553_im = _RAND_787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_554_re = _RAND_788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_554_im = _RAND_789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_555_re = _RAND_790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_555_im = _RAND_791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_556_re = _RAND_792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_556_im = _RAND_793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_557_re = _RAND_794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_557_im = _RAND_795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_558_re = _RAND_796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_558_im = _RAND_797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_559_re = _RAND_798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_559_im = _RAND_799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_560_re = _RAND_800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_560_im = _RAND_801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_561_re = _RAND_802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_561_im = _RAND_803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_562_re = _RAND_804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_562_im = _RAND_805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_563_re = _RAND_806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_563_im = _RAND_807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_564_re = _RAND_808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_564_im = _RAND_809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_565_re = _RAND_810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_565_im = _RAND_811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_566_re = _RAND_812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_566_im = _RAND_813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_567_re = _RAND_814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_567_im = _RAND_815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_568_re = _RAND_816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_568_im = _RAND_817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_569_re = _RAND_818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_569_im = _RAND_819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_570_re = _RAND_820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_570_im = _RAND_821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_571_re = _RAND_822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_571_im = _RAND_823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_572_re = _RAND_824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_572_im = _RAND_825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_573_re = _RAND_826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_573_im = _RAND_827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_574_re = _RAND_828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_574_im = _RAND_829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_575_re = _RAND_830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_575_im = _RAND_831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_576_re = _RAND_832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_576_im = _RAND_833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_577_re = _RAND_834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_577_im = _RAND_835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_578_re = _RAND_836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_578_im = _RAND_837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_579_re = _RAND_838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_579_im = _RAND_839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_580_re = _RAND_840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_580_im = _RAND_841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_581_re = _RAND_842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_581_im = _RAND_843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_582_re = _RAND_844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_582_im = _RAND_845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_583_re = _RAND_846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_583_im = _RAND_847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_584_re = _RAND_848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_584_im = _RAND_849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_585_re = _RAND_850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_585_im = _RAND_851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_586_re = _RAND_852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_586_im = _RAND_853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_587_re = _RAND_854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_587_im = _RAND_855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_588_re = _RAND_856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_588_im = _RAND_857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_589_re = _RAND_858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_589_im = _RAND_859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_590_re = _RAND_860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_590_im = _RAND_861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_591_re = _RAND_862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_591_im = _RAND_863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_592_re = _RAND_864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_592_im = _RAND_865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_593_re = _RAND_866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_593_im = _RAND_867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_594_re = _RAND_868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_594_im = _RAND_869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_595_re = _RAND_870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_595_im = _RAND_871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_596_re = _RAND_872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_596_im = _RAND_873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_597_re = _RAND_874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_597_im = _RAND_875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_598_re = _RAND_876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_598_im = _RAND_877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_599_re = _RAND_878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_599_im = _RAND_879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_600_re = _RAND_880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_600_im = _RAND_881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_601_re = _RAND_882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_601_im = _RAND_883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_602_re = _RAND_884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_602_im = _RAND_885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_603_re = _RAND_886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_603_im = _RAND_887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_604_re = _RAND_888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_604_im = _RAND_889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_605_re = _RAND_890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_605_im = _RAND_891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_606_re = _RAND_892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_606_im = _RAND_893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_607_re = _RAND_894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_607_im = _RAND_895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_608_re = _RAND_896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_608_im = _RAND_897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_609_re = _RAND_898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_609_im = _RAND_899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_610_re = _RAND_900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_610_im = _RAND_901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_611_re = _RAND_902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_611_im = _RAND_903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_612_re = _RAND_904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_612_im = _RAND_905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_613_re = _RAND_906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_613_im = _RAND_907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_614_re = _RAND_908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_614_im = _RAND_909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_615_re = _RAND_910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_615_im = _RAND_911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_616_re = _RAND_912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_616_im = _RAND_913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_617_re = _RAND_914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_617_im = _RAND_915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_618_re = _RAND_916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_618_im = _RAND_917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_619_re = _RAND_918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_619_im = _RAND_919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_620_re = _RAND_920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_620_im = _RAND_921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_621_re = _RAND_922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_621_im = _RAND_923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_622_re = _RAND_924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_622_im = _RAND_925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_623_re = _RAND_926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_623_im = _RAND_927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_624_re = _RAND_928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_624_im = _RAND_929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_625_re = _RAND_930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_625_im = _RAND_931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_626_re = _RAND_932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_626_im = _RAND_933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_627_re = _RAND_934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_627_im = _RAND_935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_628_re = _RAND_936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_628_im = _RAND_937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_629_re = _RAND_938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_629_im = _RAND_939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_630_re = _RAND_940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_630_im = _RAND_941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_631_re = _RAND_942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_631_im = _RAND_943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_632_re = _RAND_944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_632_im = _RAND_945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_633_re = _RAND_946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_633_im = _RAND_947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_634_re = _RAND_948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_634_im = _RAND_949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_635_re = _RAND_950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_635_im = _RAND_951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_636_re = _RAND_952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_636_im = _RAND_953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_637_re = _RAND_954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_637_im = _RAND_955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_638_re = _RAND_956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_638_im = _RAND_957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_639_re = _RAND_958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_639_im = _RAND_959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_640_re = _RAND_960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_640_im = _RAND_961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_641_re = _RAND_962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_641_im = _RAND_963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_642_re = _RAND_964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_642_im = _RAND_965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_643_re = _RAND_966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_643_im = _RAND_967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_644_re = _RAND_968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_644_im = _RAND_969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_645_re = _RAND_970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_645_im = _RAND_971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_646_re = _RAND_972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_646_im = _RAND_973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_647_re = _RAND_974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_647_im = _RAND_975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_648_re = _RAND_976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_648_im = _RAND_977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_649_re = _RAND_978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_649_im = _RAND_979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_650_re = _RAND_980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_650_im = _RAND_981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_651_re = _RAND_982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_651_im = _RAND_983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_652_re = _RAND_984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_652_im = _RAND_985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_653_re = _RAND_986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_653_im = _RAND_987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_654_re = _RAND_988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_654_im = _RAND_989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_655_re = _RAND_990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_655_im = _RAND_991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_656_re = _RAND_992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_656_im = _RAND_993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_657_re = _RAND_994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_657_im = _RAND_995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_658_re = _RAND_996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_658_im = _RAND_997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_659_re = _RAND_998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_659_im = _RAND_999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_660_re = _RAND_1000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_660_im = _RAND_1001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_661_re = _RAND_1002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_661_im = _RAND_1003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_662_re = _RAND_1004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_662_im = _RAND_1005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_663_re = _RAND_1006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_663_im = _RAND_1007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_664_re = _RAND_1008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_664_im = _RAND_1009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_665_re = _RAND_1010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_665_im = _RAND_1011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_666_re = _RAND_1012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_666_im = _RAND_1013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_667_re = _RAND_1014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_667_im = _RAND_1015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_668_re = _RAND_1016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_668_im = _RAND_1017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_669_re = _RAND_1018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_669_im = _RAND_1019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_670_re = _RAND_1020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_670_im = _RAND_1021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_671_re = _RAND_1022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_671_im = _RAND_1023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_672_re = _RAND_1024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_672_im = _RAND_1025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_675_re = _RAND_1026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_675_im = _RAND_1027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_676_re = _RAND_1028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_676_im = _RAND_1029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_677_re = _RAND_1030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_677_im = _RAND_1031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_678_re = _RAND_1032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_678_im = _RAND_1033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_679_re = _RAND_1034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_679_im = _RAND_1035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_680_re = _RAND_1036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_680_im = _RAND_1037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_681_re = _RAND_1038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_681_im = _RAND_1039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_682_re = _RAND_1040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_682_im = _RAND_1041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_683_re = _RAND_1042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_683_im = _RAND_1043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_684_re = _RAND_1044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_684_im = _RAND_1045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_685_re = _RAND_1046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_685_im = _RAND_1047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_686_re = _RAND_1048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_686_im = _RAND_1049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_687_re = _RAND_1050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_687_im = _RAND_1051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_688_re = _RAND_1052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_688_im = _RAND_1053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_689_re = _RAND_1054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_689_im = _RAND_1055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_690_re = _RAND_1056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_690_im = _RAND_1057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_691_re = _RAND_1058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_691_im = _RAND_1059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_692_re = _RAND_1060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_692_im = _RAND_1061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_693_re = _RAND_1062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_693_im = _RAND_1063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_694_re = _RAND_1064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_694_im = _RAND_1065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_695_re = _RAND_1066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_695_im = _RAND_1067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_696_re = _RAND_1068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_696_im = _RAND_1069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_697_re = _RAND_1070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_697_im = _RAND_1071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_698_re = _RAND_1072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_698_im = _RAND_1073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_699_re = _RAND_1074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_699_im = _RAND_1075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_700_re = _RAND_1076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_700_im = _RAND_1077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_701_re = _RAND_1078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_701_im = _RAND_1079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_702_re = _RAND_1080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_702_im = _RAND_1081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_703_re = _RAND_1082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_703_im = _RAND_1083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_704_re = _RAND_1084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_704_im = _RAND_1085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_705_re = _RAND_1086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_705_im = _RAND_1087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_706_re = _RAND_1088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_706_im = _RAND_1089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_707_re = _RAND_1090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_707_im = _RAND_1091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_708_re = _RAND_1092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_708_im = _RAND_1093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_709_re = _RAND_1094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_709_im = _RAND_1095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_710_re = _RAND_1096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_710_im = _RAND_1097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_711_re = _RAND_1098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_711_im = _RAND_1099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_712_re = _RAND_1100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_712_im = _RAND_1101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_713_re = _RAND_1102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_713_im = _RAND_1103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_714_re = _RAND_1104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_714_im = _RAND_1105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_715_re = _RAND_1106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_715_im = _RAND_1107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_716_re = _RAND_1108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_716_im = _RAND_1109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_717_re = _RAND_1110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_717_im = _RAND_1111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_718_re = _RAND_1112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_718_im = _RAND_1113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_719_re = _RAND_1114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_719_im = _RAND_1115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_720_re = _RAND_1116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_720_im = _RAND_1117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_721_re = _RAND_1118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_721_im = _RAND_1119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_722_re = _RAND_1120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_722_im = _RAND_1121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_723_re = _RAND_1122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_723_im = _RAND_1123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_724_re = _RAND_1124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_724_im = _RAND_1125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_725_re = _RAND_1126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_725_im = _RAND_1127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_726_re = _RAND_1128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_726_im = _RAND_1129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_727_re = _RAND_1130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_727_im = _RAND_1131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_728_re = _RAND_1132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_728_im = _RAND_1133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_729_re = _RAND_1134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_729_im = _RAND_1135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_730_re = _RAND_1136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_730_im = _RAND_1137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_731_re = _RAND_1138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_731_im = _RAND_1139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_732_re = _RAND_1140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_732_im = _RAND_1141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_733_re = _RAND_1142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_733_im = _RAND_1143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_734_re = _RAND_1144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_734_im = _RAND_1145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_735_re = _RAND_1146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_735_im = _RAND_1147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_736_re = _RAND_1148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_736_im = _RAND_1149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_737_re = _RAND_1150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_737_im = _RAND_1151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_738_re = _RAND_1152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_738_im = _RAND_1153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_739_re = _RAND_1154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_739_im = _RAND_1155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_740_re = _RAND_1156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_740_im = _RAND_1157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_741_re = _RAND_1158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_741_im = _RAND_1159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_742_re = _RAND_1160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_742_im = _RAND_1161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_743_re = _RAND_1162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_743_im = _RAND_1163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_744_re = _RAND_1164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_744_im = _RAND_1165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_745_re = _RAND_1166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_745_im = _RAND_1167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_746_re = _RAND_1168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_746_im = _RAND_1169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_747_re = _RAND_1170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_747_im = _RAND_1171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_748_re = _RAND_1172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_748_im = _RAND_1173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_749_re = _RAND_1174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_749_im = _RAND_1175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_750_re = _RAND_1176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_750_im = _RAND_1177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_751_re = _RAND_1178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_751_im = _RAND_1179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_752_re = _RAND_1180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_752_im = _RAND_1181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_753_re = _RAND_1182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_753_im = _RAND_1183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_754_re = _RAND_1184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_754_im = _RAND_1185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_755_re = _RAND_1186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_755_im = _RAND_1187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_756_re = _RAND_1188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_756_im = _RAND_1189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_757_re = _RAND_1190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_757_im = _RAND_1191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_758_re = _RAND_1192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_758_im = _RAND_1193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_759_re = _RAND_1194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_759_im = _RAND_1195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_760_re = _RAND_1196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_760_im = _RAND_1197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_761_re = _RAND_1198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_761_im = _RAND_1199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_762_re = _RAND_1200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_762_im = _RAND_1201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_763_re = _RAND_1202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_763_im = _RAND_1203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_764_re = _RAND_1204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_764_im = _RAND_1205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_765_re = _RAND_1206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_765_im = _RAND_1207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_766_re = _RAND_1208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_766_im = _RAND_1209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_767_re = _RAND_1210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_767_im = _RAND_1211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_768_re = _RAND_1212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_768_im = _RAND_1213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_769_re = _RAND_1214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_769_im = _RAND_1215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_770_re = _RAND_1216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_770_im = _RAND_1217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_771_re = _RAND_1218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_771_im = _RAND_1219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_772_re = _RAND_1220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_772_im = _RAND_1221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_773_re = _RAND_1222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_773_im = _RAND_1223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_774_re = _RAND_1224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_774_im = _RAND_1225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_775_re = _RAND_1226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_775_im = _RAND_1227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_776_re = _RAND_1228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_776_im = _RAND_1229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_777_re = _RAND_1230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_777_im = _RAND_1231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_778_re = _RAND_1232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_778_im = _RAND_1233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_779_re = _RAND_1234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_779_im = _RAND_1235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_780_re = _RAND_1236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_780_im = _RAND_1237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_781_re = _RAND_1238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_781_im = _RAND_1239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_782_re = _RAND_1240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_782_im = _RAND_1241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_783_re = _RAND_1242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_783_im = _RAND_1243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_784_re = _RAND_1244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_784_im = _RAND_1245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_785_re = _RAND_1246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_785_im = _RAND_1247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_786_re = _RAND_1248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_786_im = _RAND_1249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_787_re = _RAND_1250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_787_im = _RAND_1251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  _T_788_re = _RAND_1252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  _T_788_im = _RAND_1253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  _T_789_re = _RAND_1254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  _T_789_im = _RAND_1255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  _T_790_re = _RAND_1256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  _T_790_im = _RAND_1257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  _T_791_re = _RAND_1258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  _T_791_im = _RAND_1259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  _T_792_re = _RAND_1260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  _T_792_im = _RAND_1261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  _T_793_re = _RAND_1262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  _T_793_im = _RAND_1263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  _T_794_re = _RAND_1264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  _T_794_im = _RAND_1265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  _T_795_re = _RAND_1266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  _T_795_im = _RAND_1267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  _T_796_re = _RAND_1268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  _T_796_im = _RAND_1269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  _T_797_re = _RAND_1270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  _T_797_im = _RAND_1271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  _T_798_re = _RAND_1272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  _T_798_im = _RAND_1273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  _T_799_re = _RAND_1274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  _T_799_im = _RAND_1275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  _T_800_re = _RAND_1276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  _T_800_im = _RAND_1277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  _T_801_re = _RAND_1278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  _T_801_im = _RAND_1279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  _T_802_re = _RAND_1280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  _T_802_im = _RAND_1281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  _T_803_re = _RAND_1282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  _T_803_im = _RAND_1283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  _T_804_re = _RAND_1284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  _T_804_im = _RAND_1285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  _T_805_re = _RAND_1286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  _T_805_im = _RAND_1287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  _T_806_re = _RAND_1288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  _T_806_im = _RAND_1289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  _T_807_re = _RAND_1290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  _T_807_im = _RAND_1291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  _T_808_re = _RAND_1292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  _T_808_im = _RAND_1293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  _T_809_re = _RAND_1294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  _T_809_im = _RAND_1295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  _T_810_re = _RAND_1296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  _T_810_im = _RAND_1297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  _T_811_re = _RAND_1298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  _T_811_im = _RAND_1299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  _T_812_re = _RAND_1300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  _T_812_im = _RAND_1301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  _T_813_re = _RAND_1302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  _T_813_im = _RAND_1303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  _T_814_re = _RAND_1304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  _T_814_im = _RAND_1305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  _T_815_re = _RAND_1306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  _T_815_im = _RAND_1307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  _T_816_re = _RAND_1308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  _T_816_im = _RAND_1309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  _T_817_re = _RAND_1310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  _T_817_im = _RAND_1311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  _T_818_re = _RAND_1312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  _T_818_im = _RAND_1313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  _T_819_re = _RAND_1314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  _T_819_im = _RAND_1315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  _T_820_re = _RAND_1316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  _T_820_im = _RAND_1317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  _T_821_re = _RAND_1318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  _T_821_im = _RAND_1319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  _T_822_re = _RAND_1320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  _T_822_im = _RAND_1321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  _T_823_re = _RAND_1322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  _T_823_im = _RAND_1323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  _T_824_re = _RAND_1324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  _T_824_im = _RAND_1325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  _T_825_re = _RAND_1326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  _T_825_im = _RAND_1327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  _T_826_re = _RAND_1328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  _T_826_im = _RAND_1329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  _T_827_re = _RAND_1330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  _T_827_im = _RAND_1331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  _T_828_re = _RAND_1332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  _T_828_im = _RAND_1333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  _T_829_re = _RAND_1334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  _T_829_im = _RAND_1335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  _T_830_re = _RAND_1336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  _T_830_im = _RAND_1337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  _T_831_re = _RAND_1338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  _T_831_im = _RAND_1339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  _T_832_re = _RAND_1340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  _T_832_im = _RAND_1341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  _T_833_re = _RAND_1342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  _T_833_im = _RAND_1343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  _T_834_re = _RAND_1344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  _T_834_im = _RAND_1345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  _T_835_re = _RAND_1346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  _T_835_im = _RAND_1347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  _T_836_re = _RAND_1348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  _T_836_im = _RAND_1349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  _T_837_re = _RAND_1350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  _T_837_im = _RAND_1351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  _T_838_re = _RAND_1352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  _T_838_im = _RAND_1353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  _T_839_re = _RAND_1354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  _T_839_im = _RAND_1355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  _T_840_re = _RAND_1356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  _T_840_im = _RAND_1357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  _T_841_re = _RAND_1358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  _T_841_im = _RAND_1359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  _T_842_re = _RAND_1360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  _T_842_im = _RAND_1361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  _T_843_re = _RAND_1362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  _T_843_im = _RAND_1363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  _T_844_re = _RAND_1364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  _T_844_im = _RAND_1365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  _T_845_re = _RAND_1366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  _T_845_im = _RAND_1367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  _T_846_re = _RAND_1368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  _T_846_im = _RAND_1369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  _T_847_re = _RAND_1370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  _T_847_im = _RAND_1371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  _T_848_re = _RAND_1372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  _T_848_im = _RAND_1373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  _T_849_re = _RAND_1374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  _T_849_im = _RAND_1375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  _T_850_re = _RAND_1376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  _T_850_im = _RAND_1377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  _T_851_re = _RAND_1378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  _T_851_im = _RAND_1379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  _T_852_re = _RAND_1380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  _T_852_im = _RAND_1381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  _T_853_re = _RAND_1382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  _T_853_im = _RAND_1383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  _T_854_re = _RAND_1384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  _T_854_im = _RAND_1385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  _T_855_re = _RAND_1386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  _T_855_im = _RAND_1387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  _T_856_re = _RAND_1388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  _T_856_im = _RAND_1389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  _T_857_re = _RAND_1390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  _T_857_im = _RAND_1391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  _T_858_re = _RAND_1392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  _T_858_im = _RAND_1393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  _T_859_re = _RAND_1394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  _T_859_im = _RAND_1395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  _T_860_re = _RAND_1396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  _T_860_im = _RAND_1397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  _T_861_re = _RAND_1398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  _T_861_im = _RAND_1399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  _T_862_re = _RAND_1400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  _T_862_im = _RAND_1401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  _T_863_re = _RAND_1402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  _T_863_im = _RAND_1403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  _T_864_re = _RAND_1404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  _T_864_im = _RAND_1405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  _T_865_re = _RAND_1406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  _T_865_im = _RAND_1407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  _T_866_re = _RAND_1408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  _T_866_im = _RAND_1409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  _T_867_re = _RAND_1410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  _T_867_im = _RAND_1411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  _T_868_re = _RAND_1412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  _T_868_im = _RAND_1413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  _T_869_re = _RAND_1414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  _T_869_im = _RAND_1415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  _T_870_re = _RAND_1416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  _T_870_im = _RAND_1417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  _T_871_re = _RAND_1418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  _T_871_im = _RAND_1419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  _T_872_re = _RAND_1420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  _T_872_im = _RAND_1421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  _T_873_re = _RAND_1422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  _T_873_im = _RAND_1423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  _T_874_re = _RAND_1424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  _T_874_im = _RAND_1425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  _T_875_re = _RAND_1426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  _T_875_im = _RAND_1427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  _T_876_re = _RAND_1428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  _T_876_im = _RAND_1429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  _T_877_re = _RAND_1430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  _T_877_im = _RAND_1431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  _T_878_re = _RAND_1432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  _T_878_im = _RAND_1433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  _T_879_re = _RAND_1434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  _T_879_im = _RAND_1435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  _T_880_re = _RAND_1436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  _T_880_im = _RAND_1437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  _T_881_re = _RAND_1438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  _T_881_im = _RAND_1439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  _T_882_re = _RAND_1440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  _T_882_im = _RAND_1441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  _T_883_re = _RAND_1442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  _T_883_im = _RAND_1443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  _T_884_re = _RAND_1444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  _T_884_im = _RAND_1445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  _T_885_re = _RAND_1446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  _T_885_im = _RAND_1447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  _T_886_re = _RAND_1448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  _T_886_im = _RAND_1449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  _T_887_re = _RAND_1450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  _T_887_im = _RAND_1451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  _T_888_re = _RAND_1452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  _T_888_im = _RAND_1453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  _T_889_re = _RAND_1454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  _T_889_im = _RAND_1455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  _T_890_re = _RAND_1456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  _T_890_im = _RAND_1457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  _T_891_re = _RAND_1458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  _T_891_im = _RAND_1459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  _T_892_re = _RAND_1460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  _T_892_im = _RAND_1461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  _T_893_re = _RAND_1462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  _T_893_im = _RAND_1463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  _T_894_re = _RAND_1464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  _T_894_im = _RAND_1465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  _T_895_re = _RAND_1466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  _T_895_im = _RAND_1467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  _T_896_re = _RAND_1468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  _T_896_im = _RAND_1469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  _T_897_re = _RAND_1470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  _T_897_im = _RAND_1471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  _T_898_re = _RAND_1472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  _T_898_im = _RAND_1473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  _T_899_re = _RAND_1474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  _T_899_im = _RAND_1475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  _T_900_re = _RAND_1476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  _T_900_im = _RAND_1477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  _T_901_re = _RAND_1478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  _T_901_im = _RAND_1479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  _T_902_re = _RAND_1480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  _T_902_im = _RAND_1481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  _T_903_re = _RAND_1482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  _T_903_im = _RAND_1483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  _T_904_re = _RAND_1484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  _T_904_im = _RAND_1485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  _T_905_re = _RAND_1486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  _T_905_im = _RAND_1487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  _T_906_re = _RAND_1488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  _T_906_im = _RAND_1489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  _T_907_re = _RAND_1490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  _T_907_im = _RAND_1491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  _T_908_re = _RAND_1492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  _T_908_im = _RAND_1493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  _T_909_re = _RAND_1494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  _T_909_im = _RAND_1495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  _T_910_re = _RAND_1496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  _T_910_im = _RAND_1497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  _T_911_re = _RAND_1498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  _T_911_im = _RAND_1499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  _T_912_re = _RAND_1500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  _T_912_im = _RAND_1501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  _T_913_re = _RAND_1502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  _T_913_im = _RAND_1503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  _T_914_re = _RAND_1504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  _T_914_im = _RAND_1505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  _T_915_re = _RAND_1506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  _T_915_im = _RAND_1507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  _T_916_re = _RAND_1508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  _T_916_im = _RAND_1509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  _T_917_re = _RAND_1510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  _T_917_im = _RAND_1511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  _T_918_re = _RAND_1512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  _T_918_im = _RAND_1513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  _T_919_re = _RAND_1514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  _T_919_im = _RAND_1515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  _T_920_re = _RAND_1516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  _T_920_im = _RAND_1517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  _T_921_re = _RAND_1518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  _T_921_im = _RAND_1519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  _T_922_re = _RAND_1520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  _T_922_im = _RAND_1521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  _T_923_re = _RAND_1522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  _T_923_im = _RAND_1523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  _T_924_re = _RAND_1524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  _T_924_im = _RAND_1525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  _T_925_re = _RAND_1526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  _T_925_im = _RAND_1527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  _T_926_re = _RAND_1528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  _T_926_im = _RAND_1529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  _T_927_re = _RAND_1530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  _T_927_im = _RAND_1531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  _T_928_re = _RAND_1532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  _T_928_im = _RAND_1533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  _T_929_re = _RAND_1534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  _T_929_im = _RAND_1535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  _T_930_re = _RAND_1536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  _T_930_im = _RAND_1537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  _T_936_re = _RAND_1538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  _T_936_im = _RAND_1539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  _T_937_re = _RAND_1540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  _T_937_im = _RAND_1541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  _T_938_re = _RAND_1542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1543 = {1{`RANDOM}};
  _T_938_im = _RAND_1543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1544 = {1{`RANDOM}};
  _T_939_re = _RAND_1544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1545 = {1{`RANDOM}};
  _T_939_im = _RAND_1545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1546 = {1{`RANDOM}};
  _T_940_re = _RAND_1546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1547 = {1{`RANDOM}};
  _T_940_im = _RAND_1547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1548 = {1{`RANDOM}};
  _T_941_re = _RAND_1548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1549 = {1{`RANDOM}};
  _T_941_im = _RAND_1549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1550 = {1{`RANDOM}};
  _T_942_re = _RAND_1550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1551 = {1{`RANDOM}};
  _T_942_im = _RAND_1551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1552 = {1{`RANDOM}};
  _T_943_re = _RAND_1552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1553 = {1{`RANDOM}};
  _T_943_im = _RAND_1553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1554 = {1{`RANDOM}};
  _T_944_re = _RAND_1554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1555 = {1{`RANDOM}};
  _T_944_im = _RAND_1555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1556 = {1{`RANDOM}};
  _T_945_re = _RAND_1556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1557 = {1{`RANDOM}};
  _T_945_im = _RAND_1557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1558 = {1{`RANDOM}};
  _T_946_re = _RAND_1558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1559 = {1{`RANDOM}};
  _T_946_im = _RAND_1559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1560 = {1{`RANDOM}};
  _T_947_re = _RAND_1560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1561 = {1{`RANDOM}};
  _T_947_im = _RAND_1561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1562 = {1{`RANDOM}};
  _T_948_re = _RAND_1562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1563 = {1{`RANDOM}};
  _T_948_im = _RAND_1563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1564 = {1{`RANDOM}};
  _T_949_re = _RAND_1564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1565 = {1{`RANDOM}};
  _T_949_im = _RAND_1565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1566 = {1{`RANDOM}};
  _T_950_re = _RAND_1566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1567 = {1{`RANDOM}};
  _T_950_im = _RAND_1567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1568 = {1{`RANDOM}};
  _T_951_re = _RAND_1568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1569 = {1{`RANDOM}};
  _T_951_im = _RAND_1569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1570 = {1{`RANDOM}};
  _T_952_re = _RAND_1570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1571 = {1{`RANDOM}};
  _T_952_im = _RAND_1571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1572 = {1{`RANDOM}};
  _T_953_re = _RAND_1572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1573 = {1{`RANDOM}};
  _T_953_im = _RAND_1573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1574 = {1{`RANDOM}};
  _T_954_re = _RAND_1574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1575 = {1{`RANDOM}};
  _T_954_im = _RAND_1575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1576 = {1{`RANDOM}};
  _T_955_re = _RAND_1576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1577 = {1{`RANDOM}};
  _T_955_im = _RAND_1577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1578 = {1{`RANDOM}};
  _T_956_re = _RAND_1578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1579 = {1{`RANDOM}};
  _T_956_im = _RAND_1579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1580 = {1{`RANDOM}};
  _T_957_re = _RAND_1580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1581 = {1{`RANDOM}};
  _T_957_im = _RAND_1581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1582 = {1{`RANDOM}};
  _T_958_re = _RAND_1582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1583 = {1{`RANDOM}};
  _T_958_im = _RAND_1583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1584 = {1{`RANDOM}};
  _T_959_re = _RAND_1584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1585 = {1{`RANDOM}};
  _T_959_im = _RAND_1585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1586 = {1{`RANDOM}};
  _T_960_re = _RAND_1586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1587 = {1{`RANDOM}};
  _T_960_im = _RAND_1587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1588 = {1{`RANDOM}};
  _T_961_re = _RAND_1588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1589 = {1{`RANDOM}};
  _T_961_im = _RAND_1589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1590 = {1{`RANDOM}};
  _T_962_re = _RAND_1590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1591 = {1{`RANDOM}};
  _T_962_im = _RAND_1591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1592 = {1{`RANDOM}};
  _T_963_re = _RAND_1592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1593 = {1{`RANDOM}};
  _T_963_im = _RAND_1593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1594 = {1{`RANDOM}};
  _T_964_re = _RAND_1594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1595 = {1{`RANDOM}};
  _T_964_im = _RAND_1595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1596 = {1{`RANDOM}};
  _T_965_re = _RAND_1596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1597 = {1{`RANDOM}};
  _T_965_im = _RAND_1597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1598 = {1{`RANDOM}};
  _T_966_re = _RAND_1598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1599 = {1{`RANDOM}};
  _T_966_im = _RAND_1599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1600 = {1{`RANDOM}};
  _T_967_re = _RAND_1600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1601 = {1{`RANDOM}};
  _T_967_im = _RAND_1601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1602 = {1{`RANDOM}};
  _T_968_re = _RAND_1602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1603 = {1{`RANDOM}};
  _T_968_im = _RAND_1603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1604 = {1{`RANDOM}};
  _T_969_re = _RAND_1604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1605 = {1{`RANDOM}};
  _T_969_im = _RAND_1605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1606 = {1{`RANDOM}};
  _T_970_re = _RAND_1606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1607 = {1{`RANDOM}};
  _T_970_im = _RAND_1607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1608 = {1{`RANDOM}};
  _T_971_re = _RAND_1608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1609 = {1{`RANDOM}};
  _T_971_im = _RAND_1609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1610 = {1{`RANDOM}};
  _T_972_re = _RAND_1610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1611 = {1{`RANDOM}};
  _T_972_im = _RAND_1611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1612 = {1{`RANDOM}};
  _T_973_re = _RAND_1612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1613 = {1{`RANDOM}};
  _T_973_im = _RAND_1613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1614 = {1{`RANDOM}};
  _T_974_re = _RAND_1614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1615 = {1{`RANDOM}};
  _T_974_im = _RAND_1615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1616 = {1{`RANDOM}};
  _T_975_re = _RAND_1616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1617 = {1{`RANDOM}};
  _T_975_im = _RAND_1617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1618 = {1{`RANDOM}};
  _T_976_re = _RAND_1618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1619 = {1{`RANDOM}};
  _T_976_im = _RAND_1619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1620 = {1{`RANDOM}};
  _T_977_re = _RAND_1620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1621 = {1{`RANDOM}};
  _T_977_im = _RAND_1621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1622 = {1{`RANDOM}};
  _T_978_re = _RAND_1622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1623 = {1{`RANDOM}};
  _T_978_im = _RAND_1623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1624 = {1{`RANDOM}};
  _T_979_re = _RAND_1624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1625 = {1{`RANDOM}};
  _T_979_im = _RAND_1625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1626 = {1{`RANDOM}};
  _T_980_re = _RAND_1626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1627 = {1{`RANDOM}};
  _T_980_im = _RAND_1627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1628 = {1{`RANDOM}};
  _T_981_re = _RAND_1628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1629 = {1{`RANDOM}};
  _T_981_im = _RAND_1629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1630 = {1{`RANDOM}};
  _T_982_re = _RAND_1630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1631 = {1{`RANDOM}};
  _T_982_im = _RAND_1631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1632 = {1{`RANDOM}};
  _T_983_re = _RAND_1632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1633 = {1{`RANDOM}};
  _T_983_im = _RAND_1633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1634 = {1{`RANDOM}};
  _T_984_re = _RAND_1634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1635 = {1{`RANDOM}};
  _T_984_im = _RAND_1635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1636 = {1{`RANDOM}};
  _T_985_re = _RAND_1636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1637 = {1{`RANDOM}};
  _T_985_im = _RAND_1637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1638 = {1{`RANDOM}};
  _T_986_re = _RAND_1638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1639 = {1{`RANDOM}};
  _T_986_im = _RAND_1639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1640 = {1{`RANDOM}};
  _T_987_re = _RAND_1640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1641 = {1{`RANDOM}};
  _T_987_im = _RAND_1641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1642 = {1{`RANDOM}};
  _T_988_re = _RAND_1642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1643 = {1{`RANDOM}};
  _T_988_im = _RAND_1643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1644 = {1{`RANDOM}};
  _T_989_re = _RAND_1644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1645 = {1{`RANDOM}};
  _T_989_im = _RAND_1645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1646 = {1{`RANDOM}};
  _T_990_re = _RAND_1646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1647 = {1{`RANDOM}};
  _T_990_im = _RAND_1647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1648 = {1{`RANDOM}};
  _T_991_re = _RAND_1648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1649 = {1{`RANDOM}};
  _T_991_im = _RAND_1649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1650 = {1{`RANDOM}};
  _T_992_re = _RAND_1650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1651 = {1{`RANDOM}};
  _T_992_im = _RAND_1651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1652 = {1{`RANDOM}};
  _T_993_re = _RAND_1652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1653 = {1{`RANDOM}};
  _T_993_im = _RAND_1653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1654 = {1{`RANDOM}};
  _T_994_re = _RAND_1654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1655 = {1{`RANDOM}};
  _T_994_im = _RAND_1655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1656 = {1{`RANDOM}};
  _T_995_re = _RAND_1656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1657 = {1{`RANDOM}};
  _T_995_im = _RAND_1657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1658 = {1{`RANDOM}};
  _T_996_re = _RAND_1658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1659 = {1{`RANDOM}};
  _T_996_im = _RAND_1659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1660 = {1{`RANDOM}};
  _T_997_re = _RAND_1660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1661 = {1{`RANDOM}};
  _T_997_im = _RAND_1661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1662 = {1{`RANDOM}};
  _T_998_re = _RAND_1662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1663 = {1{`RANDOM}};
  _T_998_im = _RAND_1663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1664 = {1{`RANDOM}};
  _T_999_re = _RAND_1664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1665 = {1{`RANDOM}};
  _T_999_im = _RAND_1665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1666 = {1{`RANDOM}};
  _T_1000_re = _RAND_1666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1667 = {1{`RANDOM}};
  _T_1000_im = _RAND_1667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1668 = {1{`RANDOM}};
  _T_1001_re = _RAND_1668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1669 = {1{`RANDOM}};
  _T_1001_im = _RAND_1669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1670 = {1{`RANDOM}};
  _T_1002_re = _RAND_1670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1671 = {1{`RANDOM}};
  _T_1002_im = _RAND_1671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1672 = {1{`RANDOM}};
  _T_1003_re = _RAND_1672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1673 = {1{`RANDOM}};
  _T_1003_im = _RAND_1673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1674 = {1{`RANDOM}};
  _T_1004_re = _RAND_1674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1675 = {1{`RANDOM}};
  _T_1004_im = _RAND_1675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1676 = {1{`RANDOM}};
  _T_1005_re = _RAND_1676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1677 = {1{`RANDOM}};
  _T_1005_im = _RAND_1677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1678 = {1{`RANDOM}};
  _T_1006_re = _RAND_1678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1679 = {1{`RANDOM}};
  _T_1006_im = _RAND_1679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1680 = {1{`RANDOM}};
  _T_1007_re = _RAND_1680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1681 = {1{`RANDOM}};
  _T_1007_im = _RAND_1681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1682 = {1{`RANDOM}};
  _T_1008_re = _RAND_1682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1683 = {1{`RANDOM}};
  _T_1008_im = _RAND_1683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1684 = {1{`RANDOM}};
  _T_1009_re = _RAND_1684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1685 = {1{`RANDOM}};
  _T_1009_im = _RAND_1685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1686 = {1{`RANDOM}};
  _T_1010_re = _RAND_1686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1687 = {1{`RANDOM}};
  _T_1010_im = _RAND_1687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1688 = {1{`RANDOM}};
  _T_1011_re = _RAND_1688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1689 = {1{`RANDOM}};
  _T_1011_im = _RAND_1689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1690 = {1{`RANDOM}};
  _T_1012_re = _RAND_1690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1691 = {1{`RANDOM}};
  _T_1012_im = _RAND_1691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1692 = {1{`RANDOM}};
  _T_1013_re = _RAND_1692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1693 = {1{`RANDOM}};
  _T_1013_im = _RAND_1693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1694 = {1{`RANDOM}};
  _T_1014_re = _RAND_1694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1695 = {1{`RANDOM}};
  _T_1014_im = _RAND_1695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1696 = {1{`RANDOM}};
  _T_1015_re = _RAND_1696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1697 = {1{`RANDOM}};
  _T_1015_im = _RAND_1697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1698 = {1{`RANDOM}};
  _T_1016_re = _RAND_1698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1699 = {1{`RANDOM}};
  _T_1016_im = _RAND_1699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1700 = {1{`RANDOM}};
  _T_1017_re = _RAND_1700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1701 = {1{`RANDOM}};
  _T_1017_im = _RAND_1701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1702 = {1{`RANDOM}};
  _T_1018_re = _RAND_1702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1703 = {1{`RANDOM}};
  _T_1018_im = _RAND_1703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1704 = {1{`RANDOM}};
  _T_1019_re = _RAND_1704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1705 = {1{`RANDOM}};
  _T_1019_im = _RAND_1705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1706 = {1{`RANDOM}};
  _T_1020_re = _RAND_1706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1707 = {1{`RANDOM}};
  _T_1020_im = _RAND_1707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1708 = {1{`RANDOM}};
  _T_1021_re = _RAND_1708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1709 = {1{`RANDOM}};
  _T_1021_im = _RAND_1709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1710 = {1{`RANDOM}};
  _T_1022_re = _RAND_1710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1711 = {1{`RANDOM}};
  _T_1022_im = _RAND_1711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1712 = {1{`RANDOM}};
  _T_1023_re = _RAND_1712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1713 = {1{`RANDOM}};
  _T_1023_im = _RAND_1713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1714 = {1{`RANDOM}};
  _T_1024_re = _RAND_1714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1715 = {1{`RANDOM}};
  _T_1024_im = _RAND_1715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1716 = {1{`RANDOM}};
  _T_1025_re = _RAND_1716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1717 = {1{`RANDOM}};
  _T_1025_im = _RAND_1717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1718 = {1{`RANDOM}};
  _T_1026_re = _RAND_1718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1719 = {1{`RANDOM}};
  _T_1026_im = _RAND_1719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1720 = {1{`RANDOM}};
  _T_1027_re = _RAND_1720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1721 = {1{`RANDOM}};
  _T_1027_im = _RAND_1721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1722 = {1{`RANDOM}};
  _T_1028_re = _RAND_1722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1723 = {1{`RANDOM}};
  _T_1028_im = _RAND_1723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1724 = {1{`RANDOM}};
  _T_1029_re = _RAND_1724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1725 = {1{`RANDOM}};
  _T_1029_im = _RAND_1725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1726 = {1{`RANDOM}};
  _T_1030_re = _RAND_1726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1727 = {1{`RANDOM}};
  _T_1030_im = _RAND_1727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1728 = {1{`RANDOM}};
  _T_1031_re = _RAND_1728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1729 = {1{`RANDOM}};
  _T_1031_im = _RAND_1729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1730 = {1{`RANDOM}};
  _T_1032_re = _RAND_1730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1731 = {1{`RANDOM}};
  _T_1032_im = _RAND_1731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1732 = {1{`RANDOM}};
  _T_1033_re = _RAND_1732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1733 = {1{`RANDOM}};
  _T_1033_im = _RAND_1733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1734 = {1{`RANDOM}};
  _T_1034_re = _RAND_1734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1735 = {1{`RANDOM}};
  _T_1034_im = _RAND_1735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1736 = {1{`RANDOM}};
  _T_1035_re = _RAND_1736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1737 = {1{`RANDOM}};
  _T_1035_im = _RAND_1737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1738 = {1{`RANDOM}};
  _T_1036_re = _RAND_1738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1739 = {1{`RANDOM}};
  _T_1036_im = _RAND_1739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1740 = {1{`RANDOM}};
  _T_1037_re = _RAND_1740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1741 = {1{`RANDOM}};
  _T_1037_im = _RAND_1741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1742 = {1{`RANDOM}};
  _T_1038_re = _RAND_1742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1743 = {1{`RANDOM}};
  _T_1038_im = _RAND_1743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1744 = {1{`RANDOM}};
  _T_1039_re = _RAND_1744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1745 = {1{`RANDOM}};
  _T_1039_im = _RAND_1745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1746 = {1{`RANDOM}};
  _T_1040_re = _RAND_1746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1747 = {1{`RANDOM}};
  _T_1040_im = _RAND_1747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1748 = {1{`RANDOM}};
  _T_1041_re = _RAND_1748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1749 = {1{`RANDOM}};
  _T_1041_im = _RAND_1749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1750 = {1{`RANDOM}};
  _T_1042_re = _RAND_1750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1751 = {1{`RANDOM}};
  _T_1042_im = _RAND_1751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1752 = {1{`RANDOM}};
  _T_1043_re = _RAND_1752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1753 = {1{`RANDOM}};
  _T_1043_im = _RAND_1753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1754 = {1{`RANDOM}};
  _T_1044_re = _RAND_1754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1755 = {1{`RANDOM}};
  _T_1044_im = _RAND_1755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1756 = {1{`RANDOM}};
  _T_1045_re = _RAND_1756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1757 = {1{`RANDOM}};
  _T_1045_im = _RAND_1757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1758 = {1{`RANDOM}};
  _T_1046_re = _RAND_1758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1759 = {1{`RANDOM}};
  _T_1046_im = _RAND_1759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1760 = {1{`RANDOM}};
  _T_1047_re = _RAND_1760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1761 = {1{`RANDOM}};
  _T_1047_im = _RAND_1761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1762 = {1{`RANDOM}};
  _T_1048_re = _RAND_1762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1763 = {1{`RANDOM}};
  _T_1048_im = _RAND_1763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1764 = {1{`RANDOM}};
  _T_1049_re = _RAND_1764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1765 = {1{`RANDOM}};
  _T_1049_im = _RAND_1765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1766 = {1{`RANDOM}};
  _T_1050_re = _RAND_1766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1767 = {1{`RANDOM}};
  _T_1050_im = _RAND_1767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1768 = {1{`RANDOM}};
  _T_1051_re = _RAND_1768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1769 = {1{`RANDOM}};
  _T_1051_im = _RAND_1769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1770 = {1{`RANDOM}};
  _T_1052_re = _RAND_1770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1771 = {1{`RANDOM}};
  _T_1052_im = _RAND_1771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1772 = {1{`RANDOM}};
  _T_1053_re = _RAND_1772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1773 = {1{`RANDOM}};
  _T_1053_im = _RAND_1773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1774 = {1{`RANDOM}};
  _T_1054_re = _RAND_1774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1775 = {1{`RANDOM}};
  _T_1054_im = _RAND_1775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1776 = {1{`RANDOM}};
  _T_1055_re = _RAND_1776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1777 = {1{`RANDOM}};
  _T_1055_im = _RAND_1777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1778 = {1{`RANDOM}};
  _T_1056_re = _RAND_1778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1779 = {1{`RANDOM}};
  _T_1056_im = _RAND_1779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1780 = {1{`RANDOM}};
  _T_1057_re = _RAND_1780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1781 = {1{`RANDOM}};
  _T_1057_im = _RAND_1781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1782 = {1{`RANDOM}};
  _T_1058_re = _RAND_1782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1783 = {1{`RANDOM}};
  _T_1058_im = _RAND_1783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1784 = {1{`RANDOM}};
  _T_1059_re = _RAND_1784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1785 = {1{`RANDOM}};
  _T_1059_im = _RAND_1785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1786 = {1{`RANDOM}};
  _T_1060_re = _RAND_1786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1787 = {1{`RANDOM}};
  _T_1060_im = _RAND_1787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1788 = {1{`RANDOM}};
  _T_1061_re = _RAND_1788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1789 = {1{`RANDOM}};
  _T_1061_im = _RAND_1789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1790 = {1{`RANDOM}};
  _T_1062_re = _RAND_1790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1791 = {1{`RANDOM}};
  _T_1062_im = _RAND_1791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1792 = {1{`RANDOM}};
  _T_1063_re = _RAND_1792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1793 = {1{`RANDOM}};
  _T_1063_im = _RAND_1793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1794 = {1{`RANDOM}};
  _T_1064_re = _RAND_1794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1795 = {1{`RANDOM}};
  _T_1064_im = _RAND_1795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1796 = {1{`RANDOM}};
  _T_1065_re = _RAND_1796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1797 = {1{`RANDOM}};
  _T_1065_im = _RAND_1797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1798 = {1{`RANDOM}};
  _T_1066_re = _RAND_1798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1799 = {1{`RANDOM}};
  _T_1066_im = _RAND_1799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1800 = {1{`RANDOM}};
  _T_1067_re = _RAND_1800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1801 = {1{`RANDOM}};
  _T_1067_im = _RAND_1801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1802 = {1{`RANDOM}};
  _T_1068_re = _RAND_1802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1803 = {1{`RANDOM}};
  _T_1068_im = _RAND_1803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1804 = {1{`RANDOM}};
  _T_1069_re = _RAND_1804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1805 = {1{`RANDOM}};
  _T_1069_im = _RAND_1805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1806 = {1{`RANDOM}};
  _T_1070_re = _RAND_1806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1807 = {1{`RANDOM}};
  _T_1070_im = _RAND_1807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1808 = {1{`RANDOM}};
  _T_1071_re = _RAND_1808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1809 = {1{`RANDOM}};
  _T_1071_im = _RAND_1809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1810 = {1{`RANDOM}};
  _T_1072_re = _RAND_1810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1811 = {1{`RANDOM}};
  _T_1072_im = _RAND_1811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1812 = {1{`RANDOM}};
  _T_1073_re = _RAND_1812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1813 = {1{`RANDOM}};
  _T_1073_im = _RAND_1813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1814 = {1{`RANDOM}};
  _T_1074_re = _RAND_1814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1815 = {1{`RANDOM}};
  _T_1074_im = _RAND_1815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1816 = {1{`RANDOM}};
  _T_1075_re = _RAND_1816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1817 = {1{`RANDOM}};
  _T_1075_im = _RAND_1817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1818 = {1{`RANDOM}};
  _T_1076_re = _RAND_1818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1819 = {1{`RANDOM}};
  _T_1076_im = _RAND_1819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1820 = {1{`RANDOM}};
  _T_1077_re = _RAND_1820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1821 = {1{`RANDOM}};
  _T_1077_im = _RAND_1821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1822 = {1{`RANDOM}};
  _T_1078_re = _RAND_1822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1823 = {1{`RANDOM}};
  _T_1078_im = _RAND_1823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1824 = {1{`RANDOM}};
  _T_1079_re = _RAND_1824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1825 = {1{`RANDOM}};
  _T_1079_im = _RAND_1825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1826 = {1{`RANDOM}};
  _T_1080_re = _RAND_1826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1827 = {1{`RANDOM}};
  _T_1080_im = _RAND_1827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1828 = {1{`RANDOM}};
  _T_1081_re = _RAND_1828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1829 = {1{`RANDOM}};
  _T_1081_im = _RAND_1829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1830 = {1{`RANDOM}};
  _T_1082_re = _RAND_1830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1831 = {1{`RANDOM}};
  _T_1082_im = _RAND_1831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1832 = {1{`RANDOM}};
  _T_1083_re = _RAND_1832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1833 = {1{`RANDOM}};
  _T_1083_im = _RAND_1833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1834 = {1{`RANDOM}};
  _T_1084_re = _RAND_1834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1835 = {1{`RANDOM}};
  _T_1084_im = _RAND_1835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1836 = {1{`RANDOM}};
  _T_1085_re = _RAND_1836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1837 = {1{`RANDOM}};
  _T_1085_im = _RAND_1837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1838 = {1{`RANDOM}};
  _T_1086_re = _RAND_1838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1839 = {1{`RANDOM}};
  _T_1086_im = _RAND_1839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1840 = {1{`RANDOM}};
  _T_1087_re = _RAND_1840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1841 = {1{`RANDOM}};
  _T_1087_im = _RAND_1841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1842 = {1{`RANDOM}};
  _T_1088_re = _RAND_1842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1843 = {1{`RANDOM}};
  _T_1088_im = _RAND_1843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1844 = {1{`RANDOM}};
  _T_1089_re = _RAND_1844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1845 = {1{`RANDOM}};
  _T_1089_im = _RAND_1845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1846 = {1{`RANDOM}};
  _T_1090_re = _RAND_1846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1847 = {1{`RANDOM}};
  _T_1090_im = _RAND_1847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1848 = {1{`RANDOM}};
  _T_1091_re = _RAND_1848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1849 = {1{`RANDOM}};
  _T_1091_im = _RAND_1849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1850 = {1{`RANDOM}};
  _T_1092_re = _RAND_1850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1851 = {1{`RANDOM}};
  _T_1092_im = _RAND_1851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1852 = {1{`RANDOM}};
  _T_1093_re = _RAND_1852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1853 = {1{`RANDOM}};
  _T_1093_im = _RAND_1853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1854 = {1{`RANDOM}};
  _T_1094_re = _RAND_1854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1855 = {1{`RANDOM}};
  _T_1094_im = _RAND_1855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1856 = {1{`RANDOM}};
  _T_1095_re = _RAND_1856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1857 = {1{`RANDOM}};
  _T_1095_im = _RAND_1857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1858 = {1{`RANDOM}};
  _T_1096_re = _RAND_1858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1859 = {1{`RANDOM}};
  _T_1096_im = _RAND_1859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1860 = {1{`RANDOM}};
  _T_1097_re = _RAND_1860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1861 = {1{`RANDOM}};
  _T_1097_im = _RAND_1861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1862 = {1{`RANDOM}};
  _T_1098_re = _RAND_1862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1863 = {1{`RANDOM}};
  _T_1098_im = _RAND_1863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1864 = {1{`RANDOM}};
  _T_1099_re = _RAND_1864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1865 = {1{`RANDOM}};
  _T_1099_im = _RAND_1865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1866 = {1{`RANDOM}};
  _T_1100_re = _RAND_1866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1867 = {1{`RANDOM}};
  _T_1100_im = _RAND_1867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1868 = {1{`RANDOM}};
  _T_1101_re = _RAND_1868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1869 = {1{`RANDOM}};
  _T_1101_im = _RAND_1869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1870 = {1{`RANDOM}};
  _T_1102_re = _RAND_1870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1871 = {1{`RANDOM}};
  _T_1102_im = _RAND_1871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1872 = {1{`RANDOM}};
  _T_1103_re = _RAND_1872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1873 = {1{`RANDOM}};
  _T_1103_im = _RAND_1873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1874 = {1{`RANDOM}};
  _T_1104_re = _RAND_1874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1875 = {1{`RANDOM}};
  _T_1104_im = _RAND_1875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1876 = {1{`RANDOM}};
  _T_1105_re = _RAND_1876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1877 = {1{`RANDOM}};
  _T_1105_im = _RAND_1877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1878 = {1{`RANDOM}};
  _T_1106_re = _RAND_1878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1879 = {1{`RANDOM}};
  _T_1106_im = _RAND_1879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1880 = {1{`RANDOM}};
  _T_1107_re = _RAND_1880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1881 = {1{`RANDOM}};
  _T_1107_im = _RAND_1881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1882 = {1{`RANDOM}};
  _T_1108_re = _RAND_1882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1883 = {1{`RANDOM}};
  _T_1108_im = _RAND_1883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1884 = {1{`RANDOM}};
  _T_1109_re = _RAND_1884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1885 = {1{`RANDOM}};
  _T_1109_im = _RAND_1885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1886 = {1{`RANDOM}};
  _T_1110_re = _RAND_1886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1887 = {1{`RANDOM}};
  _T_1110_im = _RAND_1887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1888 = {1{`RANDOM}};
  _T_1111_re = _RAND_1888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1889 = {1{`RANDOM}};
  _T_1111_im = _RAND_1889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1890 = {1{`RANDOM}};
  _T_1112_re = _RAND_1890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1891 = {1{`RANDOM}};
  _T_1112_im = _RAND_1891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1892 = {1{`RANDOM}};
  _T_1113_re = _RAND_1892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1893 = {1{`RANDOM}};
  _T_1113_im = _RAND_1893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1894 = {1{`RANDOM}};
  _T_1114_re = _RAND_1894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1895 = {1{`RANDOM}};
  _T_1114_im = _RAND_1895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1896 = {1{`RANDOM}};
  _T_1115_re = _RAND_1896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1897 = {1{`RANDOM}};
  _T_1115_im = _RAND_1897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1898 = {1{`RANDOM}};
  _T_1116_re = _RAND_1898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1899 = {1{`RANDOM}};
  _T_1116_im = _RAND_1899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1900 = {1{`RANDOM}};
  _T_1117_re = _RAND_1900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1901 = {1{`RANDOM}};
  _T_1117_im = _RAND_1901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1902 = {1{`RANDOM}};
  _T_1118_re = _RAND_1902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1903 = {1{`RANDOM}};
  _T_1118_im = _RAND_1903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1904 = {1{`RANDOM}};
  _T_1119_re = _RAND_1904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1905 = {1{`RANDOM}};
  _T_1119_im = _RAND_1905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1906 = {1{`RANDOM}};
  _T_1120_re = _RAND_1906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1907 = {1{`RANDOM}};
  _T_1120_im = _RAND_1907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1908 = {1{`RANDOM}};
  _T_1121_re = _RAND_1908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1909 = {1{`RANDOM}};
  _T_1121_im = _RAND_1909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1910 = {1{`RANDOM}};
  _T_1122_re = _RAND_1910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1911 = {1{`RANDOM}};
  _T_1122_im = _RAND_1911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1912 = {1{`RANDOM}};
  _T_1123_re = _RAND_1912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1913 = {1{`RANDOM}};
  _T_1123_im = _RAND_1913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1914 = {1{`RANDOM}};
  _T_1124_re = _RAND_1914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1915 = {1{`RANDOM}};
  _T_1124_im = _RAND_1915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1916 = {1{`RANDOM}};
  _T_1125_re = _RAND_1916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1917 = {1{`RANDOM}};
  _T_1125_im = _RAND_1917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1918 = {1{`RANDOM}};
  _T_1126_re = _RAND_1918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1919 = {1{`RANDOM}};
  _T_1126_im = _RAND_1919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1920 = {1{`RANDOM}};
  _T_1127_re = _RAND_1920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1921 = {1{`RANDOM}};
  _T_1127_im = _RAND_1921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1922 = {1{`RANDOM}};
  _T_1128_re = _RAND_1922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1923 = {1{`RANDOM}};
  _T_1128_im = _RAND_1923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1924 = {1{`RANDOM}};
  _T_1129_re = _RAND_1924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1925 = {1{`RANDOM}};
  _T_1129_im = _RAND_1925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1926 = {1{`RANDOM}};
  _T_1130_re = _RAND_1926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1927 = {1{`RANDOM}};
  _T_1130_im = _RAND_1927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1928 = {1{`RANDOM}};
  _T_1131_re = _RAND_1928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1929 = {1{`RANDOM}};
  _T_1131_im = _RAND_1929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1930 = {1{`RANDOM}};
  _T_1132_re = _RAND_1930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1931 = {1{`RANDOM}};
  _T_1132_im = _RAND_1931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1932 = {1{`RANDOM}};
  _T_1133_re = _RAND_1932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1933 = {1{`RANDOM}};
  _T_1133_im = _RAND_1933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1934 = {1{`RANDOM}};
  _T_1134_re = _RAND_1934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1935 = {1{`RANDOM}};
  _T_1134_im = _RAND_1935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1936 = {1{`RANDOM}};
  _T_1135_re = _RAND_1936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1937 = {1{`RANDOM}};
  _T_1135_im = _RAND_1937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1938 = {1{`RANDOM}};
  _T_1136_re = _RAND_1938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1939 = {1{`RANDOM}};
  _T_1136_im = _RAND_1939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1940 = {1{`RANDOM}};
  _T_1137_re = _RAND_1940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1941 = {1{`RANDOM}};
  _T_1137_im = _RAND_1941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1942 = {1{`RANDOM}};
  _T_1138_re = _RAND_1942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1943 = {1{`RANDOM}};
  _T_1138_im = _RAND_1943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1944 = {1{`RANDOM}};
  _T_1139_re = _RAND_1944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1945 = {1{`RANDOM}};
  _T_1139_im = _RAND_1945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1946 = {1{`RANDOM}};
  _T_1140_re = _RAND_1946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1947 = {1{`RANDOM}};
  _T_1140_im = _RAND_1947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1948 = {1{`RANDOM}};
  _T_1141_re = _RAND_1948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1949 = {1{`RANDOM}};
  _T_1141_im = _RAND_1949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1950 = {1{`RANDOM}};
  _T_1142_re = _RAND_1950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1951 = {1{`RANDOM}};
  _T_1142_im = _RAND_1951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1952 = {1{`RANDOM}};
  _T_1143_re = _RAND_1952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1953 = {1{`RANDOM}};
  _T_1143_im = _RAND_1953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1954 = {1{`RANDOM}};
  _T_1144_re = _RAND_1954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1955 = {1{`RANDOM}};
  _T_1144_im = _RAND_1955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1956 = {1{`RANDOM}};
  _T_1145_re = _RAND_1956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1957 = {1{`RANDOM}};
  _T_1145_im = _RAND_1957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1958 = {1{`RANDOM}};
  _T_1146_re = _RAND_1958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1959 = {1{`RANDOM}};
  _T_1146_im = _RAND_1959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1960 = {1{`RANDOM}};
  _T_1147_re = _RAND_1960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1961 = {1{`RANDOM}};
  _T_1147_im = _RAND_1961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1962 = {1{`RANDOM}};
  _T_1148_re = _RAND_1962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1963 = {1{`RANDOM}};
  _T_1148_im = _RAND_1963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1964 = {1{`RANDOM}};
  _T_1149_re = _RAND_1964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1965 = {1{`RANDOM}};
  _T_1149_im = _RAND_1965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1966 = {1{`RANDOM}};
  _T_1150_re = _RAND_1966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1967 = {1{`RANDOM}};
  _T_1150_im = _RAND_1967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1968 = {1{`RANDOM}};
  _T_1151_re = _RAND_1968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1969 = {1{`RANDOM}};
  _T_1151_im = _RAND_1969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1970 = {1{`RANDOM}};
  _T_1152_re = _RAND_1970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1971 = {1{`RANDOM}};
  _T_1152_im = _RAND_1971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1972 = {1{`RANDOM}};
  _T_1153_re = _RAND_1972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1973 = {1{`RANDOM}};
  _T_1153_im = _RAND_1973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1974 = {1{`RANDOM}};
  _T_1154_re = _RAND_1974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1975 = {1{`RANDOM}};
  _T_1154_im = _RAND_1975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1976 = {1{`RANDOM}};
  _T_1155_re = _RAND_1976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1977 = {1{`RANDOM}};
  _T_1155_im = _RAND_1977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1978 = {1{`RANDOM}};
  _T_1156_re = _RAND_1978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1979 = {1{`RANDOM}};
  _T_1156_im = _RAND_1979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1980 = {1{`RANDOM}};
  _T_1157_re = _RAND_1980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1981 = {1{`RANDOM}};
  _T_1157_im = _RAND_1981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1982 = {1{`RANDOM}};
  _T_1158_re = _RAND_1982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1983 = {1{`RANDOM}};
  _T_1158_im = _RAND_1983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1984 = {1{`RANDOM}};
  _T_1159_re = _RAND_1984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1985 = {1{`RANDOM}};
  _T_1159_im = _RAND_1985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1986 = {1{`RANDOM}};
  _T_1160_re = _RAND_1986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1987 = {1{`RANDOM}};
  _T_1160_im = _RAND_1987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1988 = {1{`RANDOM}};
  _T_1161_re = _RAND_1988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1989 = {1{`RANDOM}};
  _T_1161_im = _RAND_1989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1990 = {1{`RANDOM}};
  _T_1162_re = _RAND_1990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1991 = {1{`RANDOM}};
  _T_1162_im = _RAND_1991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1992 = {1{`RANDOM}};
  _T_1163_re = _RAND_1992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1993 = {1{`RANDOM}};
  _T_1163_im = _RAND_1993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1994 = {1{`RANDOM}};
  _T_1164_re = _RAND_1994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1995 = {1{`RANDOM}};
  _T_1164_im = _RAND_1995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1996 = {1{`RANDOM}};
  _T_1165_re = _RAND_1996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1997 = {1{`RANDOM}};
  _T_1165_im = _RAND_1997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1998 = {1{`RANDOM}};
  _T_1166_re = _RAND_1998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1999 = {1{`RANDOM}};
  _T_1166_im = _RAND_1999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2000 = {1{`RANDOM}};
  _T_1167_re = _RAND_2000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2001 = {1{`RANDOM}};
  _T_1167_im = _RAND_2001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2002 = {1{`RANDOM}};
  _T_1168_re = _RAND_2002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2003 = {1{`RANDOM}};
  _T_1168_im = _RAND_2003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2004 = {1{`RANDOM}};
  _T_1169_re = _RAND_2004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2005 = {1{`RANDOM}};
  _T_1169_im = _RAND_2005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2006 = {1{`RANDOM}};
  _T_1170_re = _RAND_2006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2007 = {1{`RANDOM}};
  _T_1170_im = _RAND_2007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2008 = {1{`RANDOM}};
  _T_1171_re = _RAND_2008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2009 = {1{`RANDOM}};
  _T_1171_im = _RAND_2009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2010 = {1{`RANDOM}};
  _T_1172_re = _RAND_2010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2011 = {1{`RANDOM}};
  _T_1172_im = _RAND_2011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2012 = {1{`RANDOM}};
  _T_1173_re = _RAND_2012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2013 = {1{`RANDOM}};
  _T_1173_im = _RAND_2013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2014 = {1{`RANDOM}};
  _T_1174_re = _RAND_2014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2015 = {1{`RANDOM}};
  _T_1174_im = _RAND_2015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2016 = {1{`RANDOM}};
  _T_1175_re = _RAND_2016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2017 = {1{`RANDOM}};
  _T_1175_im = _RAND_2017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2018 = {1{`RANDOM}};
  _T_1176_re = _RAND_2018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2019 = {1{`RANDOM}};
  _T_1176_im = _RAND_2019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2020 = {1{`RANDOM}};
  _T_1177_re = _RAND_2020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2021 = {1{`RANDOM}};
  _T_1177_im = _RAND_2021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2022 = {1{`RANDOM}};
  _T_1178_re = _RAND_2022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2023 = {1{`RANDOM}};
  _T_1178_im = _RAND_2023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2024 = {1{`RANDOM}};
  _T_1179_re = _RAND_2024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2025 = {1{`RANDOM}};
  _T_1179_im = _RAND_2025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2026 = {1{`RANDOM}};
  _T_1180_re = _RAND_2026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2027 = {1{`RANDOM}};
  _T_1180_im = _RAND_2027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2028 = {1{`RANDOM}};
  _T_1181_re = _RAND_2028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2029 = {1{`RANDOM}};
  _T_1181_im = _RAND_2029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2030 = {1{`RANDOM}};
  _T_1182_re = _RAND_2030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2031 = {1{`RANDOM}};
  _T_1182_im = _RAND_2031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2032 = {1{`RANDOM}};
  _T_1183_re = _RAND_2032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2033 = {1{`RANDOM}};
  _T_1183_im = _RAND_2033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2034 = {1{`RANDOM}};
  _T_1184_re = _RAND_2034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2035 = {1{`RANDOM}};
  _T_1184_im = _RAND_2035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2036 = {1{`RANDOM}};
  _T_1185_re = _RAND_2036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2037 = {1{`RANDOM}};
  _T_1185_im = _RAND_2037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2038 = {1{`RANDOM}};
  _T_1186_re = _RAND_2038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2039 = {1{`RANDOM}};
  _T_1186_im = _RAND_2039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2040 = {1{`RANDOM}};
  _T_1187_re = _RAND_2040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2041 = {1{`RANDOM}};
  _T_1187_im = _RAND_2041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2042 = {1{`RANDOM}};
  _T_1188_re = _RAND_2042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2043 = {1{`RANDOM}};
  _T_1188_im = _RAND_2043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2044 = {1{`RANDOM}};
  _T_1189_re = _RAND_2044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2045 = {1{`RANDOM}};
  _T_1189_im = _RAND_2045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2046 = {1{`RANDOM}};
  _T_1190_re = _RAND_2046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2047 = {1{`RANDOM}};
  _T_1190_im = _RAND_2047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2048 = {1{`RANDOM}};
  _T_1191_re = _RAND_2048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2049 = {1{`RANDOM}};
  _T_1191_im = _RAND_2049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2050 = {1{`RANDOM}};
  _T_1194_re = _RAND_2050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2051 = {1{`RANDOM}};
  _T_1194_im = _RAND_2051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2052 = {1{`RANDOM}};
  _T_1195_re = _RAND_2052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2053 = {1{`RANDOM}};
  _T_1195_im = _RAND_2053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2054 = {1{`RANDOM}};
  _T_1196_re = _RAND_2054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2055 = {1{`RANDOM}};
  _T_1196_im = _RAND_2055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2056 = {1{`RANDOM}};
  _T_1197_re = _RAND_2056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2057 = {1{`RANDOM}};
  _T_1197_im = _RAND_2057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2058 = {1{`RANDOM}};
  _T_1198_re = _RAND_2058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2059 = {1{`RANDOM}};
  _T_1198_im = _RAND_2059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2060 = {1{`RANDOM}};
  _T_1199_re = _RAND_2060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2061 = {1{`RANDOM}};
  _T_1199_im = _RAND_2061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2062 = {1{`RANDOM}};
  _T_1200_re = _RAND_2062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2063 = {1{`RANDOM}};
  _T_1200_im = _RAND_2063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2064 = {1{`RANDOM}};
  _T_1201_re = _RAND_2064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2065 = {1{`RANDOM}};
  _T_1201_im = _RAND_2065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2066 = {1{`RANDOM}};
  _T_1202_re = _RAND_2066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2067 = {1{`RANDOM}};
  _T_1202_im = _RAND_2067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2068 = {1{`RANDOM}};
  _T_1203_re = _RAND_2068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2069 = {1{`RANDOM}};
  _T_1203_im = _RAND_2069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2070 = {1{`RANDOM}};
  _T_1204_re = _RAND_2070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2071 = {1{`RANDOM}};
  _T_1204_im = _RAND_2071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2072 = {1{`RANDOM}};
  _T_1205_re = _RAND_2072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2073 = {1{`RANDOM}};
  _T_1205_im = _RAND_2073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2074 = {1{`RANDOM}};
  _T_1206_re = _RAND_2074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2075 = {1{`RANDOM}};
  _T_1206_im = _RAND_2075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2076 = {1{`RANDOM}};
  _T_1207_re = _RAND_2076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2077 = {1{`RANDOM}};
  _T_1207_im = _RAND_2077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2078 = {1{`RANDOM}};
  _T_1208_re = _RAND_2078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2079 = {1{`RANDOM}};
  _T_1208_im = _RAND_2079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2080 = {1{`RANDOM}};
  _T_1209_re = _RAND_2080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2081 = {1{`RANDOM}};
  _T_1209_im = _RAND_2081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2082 = {1{`RANDOM}};
  _T_1210_re = _RAND_2082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2083 = {1{`RANDOM}};
  _T_1210_im = _RAND_2083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2084 = {1{`RANDOM}};
  _T_1211_re = _RAND_2084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2085 = {1{`RANDOM}};
  _T_1211_im = _RAND_2085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2086 = {1{`RANDOM}};
  _T_1212_re = _RAND_2086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2087 = {1{`RANDOM}};
  _T_1212_im = _RAND_2087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2088 = {1{`RANDOM}};
  _T_1213_re = _RAND_2088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2089 = {1{`RANDOM}};
  _T_1213_im = _RAND_2089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2090 = {1{`RANDOM}};
  _T_1214_re = _RAND_2090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2091 = {1{`RANDOM}};
  _T_1214_im = _RAND_2091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2092 = {1{`RANDOM}};
  _T_1215_re = _RAND_2092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2093 = {1{`RANDOM}};
  _T_1215_im = _RAND_2093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2094 = {1{`RANDOM}};
  _T_1216_re = _RAND_2094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2095 = {1{`RANDOM}};
  _T_1216_im = _RAND_2095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2096 = {1{`RANDOM}};
  _T_1217_re = _RAND_2096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2097 = {1{`RANDOM}};
  _T_1217_im = _RAND_2097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2098 = {1{`RANDOM}};
  _T_1218_re = _RAND_2098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2099 = {1{`RANDOM}};
  _T_1218_im = _RAND_2099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2100 = {1{`RANDOM}};
  _T_1219_re = _RAND_2100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2101 = {1{`RANDOM}};
  _T_1219_im = _RAND_2101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2102 = {1{`RANDOM}};
  _T_1220_re = _RAND_2102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2103 = {1{`RANDOM}};
  _T_1220_im = _RAND_2103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2104 = {1{`RANDOM}};
  _T_1221_re = _RAND_2104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2105 = {1{`RANDOM}};
  _T_1221_im = _RAND_2105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2106 = {1{`RANDOM}};
  _T_1222_re = _RAND_2106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2107 = {1{`RANDOM}};
  _T_1222_im = _RAND_2107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2108 = {1{`RANDOM}};
  _T_1223_re = _RAND_2108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2109 = {1{`RANDOM}};
  _T_1223_im = _RAND_2109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2110 = {1{`RANDOM}};
  _T_1224_re = _RAND_2110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2111 = {1{`RANDOM}};
  _T_1224_im = _RAND_2111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2112 = {1{`RANDOM}};
  _T_1225_re = _RAND_2112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2113 = {1{`RANDOM}};
  _T_1225_im = _RAND_2113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2114 = {1{`RANDOM}};
  _T_1226_re = _RAND_2114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2115 = {1{`RANDOM}};
  _T_1226_im = _RAND_2115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2116 = {1{`RANDOM}};
  _T_1227_re = _RAND_2116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2117 = {1{`RANDOM}};
  _T_1227_im = _RAND_2117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2118 = {1{`RANDOM}};
  _T_1228_re = _RAND_2118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2119 = {1{`RANDOM}};
  _T_1228_im = _RAND_2119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2120 = {1{`RANDOM}};
  _T_1229_re = _RAND_2120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2121 = {1{`RANDOM}};
  _T_1229_im = _RAND_2121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2122 = {1{`RANDOM}};
  _T_1230_re = _RAND_2122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2123 = {1{`RANDOM}};
  _T_1230_im = _RAND_2123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2124 = {1{`RANDOM}};
  _T_1231_re = _RAND_2124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2125 = {1{`RANDOM}};
  _T_1231_im = _RAND_2125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2126 = {1{`RANDOM}};
  _T_1232_re = _RAND_2126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2127 = {1{`RANDOM}};
  _T_1232_im = _RAND_2127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2128 = {1{`RANDOM}};
  _T_1233_re = _RAND_2128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2129 = {1{`RANDOM}};
  _T_1233_im = _RAND_2129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2130 = {1{`RANDOM}};
  _T_1234_re = _RAND_2130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2131 = {1{`RANDOM}};
  _T_1234_im = _RAND_2131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2132 = {1{`RANDOM}};
  _T_1235_re = _RAND_2132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2133 = {1{`RANDOM}};
  _T_1235_im = _RAND_2133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2134 = {1{`RANDOM}};
  _T_1236_re = _RAND_2134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2135 = {1{`RANDOM}};
  _T_1236_im = _RAND_2135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2136 = {1{`RANDOM}};
  _T_1237_re = _RAND_2136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2137 = {1{`RANDOM}};
  _T_1237_im = _RAND_2137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2138 = {1{`RANDOM}};
  _T_1238_re = _RAND_2138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2139 = {1{`RANDOM}};
  _T_1238_im = _RAND_2139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2140 = {1{`RANDOM}};
  _T_1239_re = _RAND_2140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2141 = {1{`RANDOM}};
  _T_1239_im = _RAND_2141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2142 = {1{`RANDOM}};
  _T_1240_re = _RAND_2142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2143 = {1{`RANDOM}};
  _T_1240_im = _RAND_2143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2144 = {1{`RANDOM}};
  _T_1241_re = _RAND_2144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2145 = {1{`RANDOM}};
  _T_1241_im = _RAND_2145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2146 = {1{`RANDOM}};
  _T_1242_re = _RAND_2146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2147 = {1{`RANDOM}};
  _T_1242_im = _RAND_2147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2148 = {1{`RANDOM}};
  _T_1243_re = _RAND_2148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2149 = {1{`RANDOM}};
  _T_1243_im = _RAND_2149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2150 = {1{`RANDOM}};
  _T_1244_re = _RAND_2150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2151 = {1{`RANDOM}};
  _T_1244_im = _RAND_2151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2152 = {1{`RANDOM}};
  _T_1245_re = _RAND_2152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2153 = {1{`RANDOM}};
  _T_1245_im = _RAND_2153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2154 = {1{`RANDOM}};
  _T_1246_re = _RAND_2154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2155 = {1{`RANDOM}};
  _T_1246_im = _RAND_2155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2156 = {1{`RANDOM}};
  _T_1247_re = _RAND_2156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2157 = {1{`RANDOM}};
  _T_1247_im = _RAND_2157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2158 = {1{`RANDOM}};
  _T_1248_re = _RAND_2158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2159 = {1{`RANDOM}};
  _T_1248_im = _RAND_2159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2160 = {1{`RANDOM}};
  _T_1249_re = _RAND_2160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2161 = {1{`RANDOM}};
  _T_1249_im = _RAND_2161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2162 = {1{`RANDOM}};
  _T_1250_re = _RAND_2162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2163 = {1{`RANDOM}};
  _T_1250_im = _RAND_2163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2164 = {1{`RANDOM}};
  _T_1251_re = _RAND_2164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2165 = {1{`RANDOM}};
  _T_1251_im = _RAND_2165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2166 = {1{`RANDOM}};
  _T_1252_re = _RAND_2166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2167 = {1{`RANDOM}};
  _T_1252_im = _RAND_2167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2168 = {1{`RANDOM}};
  _T_1253_re = _RAND_2168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2169 = {1{`RANDOM}};
  _T_1253_im = _RAND_2169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2170 = {1{`RANDOM}};
  _T_1254_re = _RAND_2170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2171 = {1{`RANDOM}};
  _T_1254_im = _RAND_2171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2172 = {1{`RANDOM}};
  _T_1255_re = _RAND_2172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2173 = {1{`RANDOM}};
  _T_1255_im = _RAND_2173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2174 = {1{`RANDOM}};
  _T_1256_re = _RAND_2174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2175 = {1{`RANDOM}};
  _T_1256_im = _RAND_2175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2176 = {1{`RANDOM}};
  _T_1257_re = _RAND_2176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2177 = {1{`RANDOM}};
  _T_1257_im = _RAND_2177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2178 = {1{`RANDOM}};
  _T_1258_re = _RAND_2178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2179 = {1{`RANDOM}};
  _T_1258_im = _RAND_2179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2180 = {1{`RANDOM}};
  _T_1259_re = _RAND_2180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2181 = {1{`RANDOM}};
  _T_1259_im = _RAND_2181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2182 = {1{`RANDOM}};
  _T_1260_re = _RAND_2182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2183 = {1{`RANDOM}};
  _T_1260_im = _RAND_2183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2184 = {1{`RANDOM}};
  _T_1261_re = _RAND_2184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2185 = {1{`RANDOM}};
  _T_1261_im = _RAND_2185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2186 = {1{`RANDOM}};
  _T_1262_re = _RAND_2186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2187 = {1{`RANDOM}};
  _T_1262_im = _RAND_2187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2188 = {1{`RANDOM}};
  _T_1263_re = _RAND_2188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2189 = {1{`RANDOM}};
  _T_1263_im = _RAND_2189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2190 = {1{`RANDOM}};
  _T_1264_re = _RAND_2190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2191 = {1{`RANDOM}};
  _T_1264_im = _RAND_2191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2192 = {1{`RANDOM}};
  _T_1265_re = _RAND_2192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2193 = {1{`RANDOM}};
  _T_1265_im = _RAND_2193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2194 = {1{`RANDOM}};
  _T_1266_re = _RAND_2194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2195 = {1{`RANDOM}};
  _T_1266_im = _RAND_2195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2196 = {1{`RANDOM}};
  _T_1267_re = _RAND_2196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2197 = {1{`RANDOM}};
  _T_1267_im = _RAND_2197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2198 = {1{`RANDOM}};
  _T_1268_re = _RAND_2198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2199 = {1{`RANDOM}};
  _T_1268_im = _RAND_2199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2200 = {1{`RANDOM}};
  _T_1269_re = _RAND_2200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2201 = {1{`RANDOM}};
  _T_1269_im = _RAND_2201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2202 = {1{`RANDOM}};
  _T_1270_re = _RAND_2202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2203 = {1{`RANDOM}};
  _T_1270_im = _RAND_2203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2204 = {1{`RANDOM}};
  _T_1271_re = _RAND_2204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2205 = {1{`RANDOM}};
  _T_1271_im = _RAND_2205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2206 = {1{`RANDOM}};
  _T_1272_re = _RAND_2206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2207 = {1{`RANDOM}};
  _T_1272_im = _RAND_2207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2208 = {1{`RANDOM}};
  _T_1273_re = _RAND_2208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2209 = {1{`RANDOM}};
  _T_1273_im = _RAND_2209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2210 = {1{`RANDOM}};
  _T_1274_re = _RAND_2210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2211 = {1{`RANDOM}};
  _T_1274_im = _RAND_2211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2212 = {1{`RANDOM}};
  _T_1275_re = _RAND_2212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2213 = {1{`RANDOM}};
  _T_1275_im = _RAND_2213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2214 = {1{`RANDOM}};
  _T_1276_re = _RAND_2214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2215 = {1{`RANDOM}};
  _T_1276_im = _RAND_2215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2216 = {1{`RANDOM}};
  _T_1277_re = _RAND_2216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2217 = {1{`RANDOM}};
  _T_1277_im = _RAND_2217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2218 = {1{`RANDOM}};
  _T_1278_re = _RAND_2218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2219 = {1{`RANDOM}};
  _T_1278_im = _RAND_2219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2220 = {1{`RANDOM}};
  _T_1279_re = _RAND_2220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2221 = {1{`RANDOM}};
  _T_1279_im = _RAND_2221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2222 = {1{`RANDOM}};
  _T_1280_re = _RAND_2222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2223 = {1{`RANDOM}};
  _T_1280_im = _RAND_2223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2224 = {1{`RANDOM}};
  _T_1281_re = _RAND_2224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2225 = {1{`RANDOM}};
  _T_1281_im = _RAND_2225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2226 = {1{`RANDOM}};
  _T_1282_re = _RAND_2226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2227 = {1{`RANDOM}};
  _T_1282_im = _RAND_2227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2228 = {1{`RANDOM}};
  _T_1283_re = _RAND_2228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2229 = {1{`RANDOM}};
  _T_1283_im = _RAND_2229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2230 = {1{`RANDOM}};
  _T_1284_re = _RAND_2230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2231 = {1{`RANDOM}};
  _T_1284_im = _RAND_2231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2232 = {1{`RANDOM}};
  _T_1285_re = _RAND_2232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2233 = {1{`RANDOM}};
  _T_1285_im = _RAND_2233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2234 = {1{`RANDOM}};
  _T_1286_re = _RAND_2234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2235 = {1{`RANDOM}};
  _T_1286_im = _RAND_2235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2236 = {1{`RANDOM}};
  _T_1287_re = _RAND_2236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2237 = {1{`RANDOM}};
  _T_1287_im = _RAND_2237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2238 = {1{`RANDOM}};
  _T_1288_re = _RAND_2238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2239 = {1{`RANDOM}};
  _T_1288_im = _RAND_2239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2240 = {1{`RANDOM}};
  _T_1289_re = _RAND_2240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2241 = {1{`RANDOM}};
  _T_1289_im = _RAND_2241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2242 = {1{`RANDOM}};
  _T_1290_re = _RAND_2242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2243 = {1{`RANDOM}};
  _T_1290_im = _RAND_2243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2244 = {1{`RANDOM}};
  _T_1291_re = _RAND_2244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2245 = {1{`RANDOM}};
  _T_1291_im = _RAND_2245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2246 = {1{`RANDOM}};
  _T_1292_re = _RAND_2246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2247 = {1{`RANDOM}};
  _T_1292_im = _RAND_2247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2248 = {1{`RANDOM}};
  _T_1293_re = _RAND_2248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2249 = {1{`RANDOM}};
  _T_1293_im = _RAND_2249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2250 = {1{`RANDOM}};
  _T_1294_re = _RAND_2250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2251 = {1{`RANDOM}};
  _T_1294_im = _RAND_2251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2252 = {1{`RANDOM}};
  _T_1295_re = _RAND_2252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2253 = {1{`RANDOM}};
  _T_1295_im = _RAND_2253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2254 = {1{`RANDOM}};
  _T_1296_re = _RAND_2254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2255 = {1{`RANDOM}};
  _T_1296_im = _RAND_2255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2256 = {1{`RANDOM}};
  _T_1297_re = _RAND_2256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2257 = {1{`RANDOM}};
  _T_1297_im = _RAND_2257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2258 = {1{`RANDOM}};
  _T_1298_re = _RAND_2258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2259 = {1{`RANDOM}};
  _T_1298_im = _RAND_2259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2260 = {1{`RANDOM}};
  _T_1299_re = _RAND_2260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2261 = {1{`RANDOM}};
  _T_1299_im = _RAND_2261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2262 = {1{`RANDOM}};
  _T_1300_re = _RAND_2262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2263 = {1{`RANDOM}};
  _T_1300_im = _RAND_2263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2264 = {1{`RANDOM}};
  _T_1301_re = _RAND_2264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2265 = {1{`RANDOM}};
  _T_1301_im = _RAND_2265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2266 = {1{`RANDOM}};
  _T_1302_re = _RAND_2266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2267 = {1{`RANDOM}};
  _T_1302_im = _RAND_2267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2268 = {1{`RANDOM}};
  _T_1303_re = _RAND_2268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2269 = {1{`RANDOM}};
  _T_1303_im = _RAND_2269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2270 = {1{`RANDOM}};
  _T_1304_re = _RAND_2270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2271 = {1{`RANDOM}};
  _T_1304_im = _RAND_2271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2272 = {1{`RANDOM}};
  _T_1305_re = _RAND_2272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2273 = {1{`RANDOM}};
  _T_1305_im = _RAND_2273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2274 = {1{`RANDOM}};
  _T_1306_re = _RAND_2274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2275 = {1{`RANDOM}};
  _T_1306_im = _RAND_2275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2276 = {1{`RANDOM}};
  _T_1307_re = _RAND_2276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2277 = {1{`RANDOM}};
  _T_1307_im = _RAND_2277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2278 = {1{`RANDOM}};
  _T_1308_re = _RAND_2278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2279 = {1{`RANDOM}};
  _T_1308_im = _RAND_2279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2280 = {1{`RANDOM}};
  _T_1309_re = _RAND_2280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2281 = {1{`RANDOM}};
  _T_1309_im = _RAND_2281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2282 = {1{`RANDOM}};
  _T_1310_re = _RAND_2282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2283 = {1{`RANDOM}};
  _T_1310_im = _RAND_2283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2284 = {1{`RANDOM}};
  _T_1311_re = _RAND_2284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2285 = {1{`RANDOM}};
  _T_1311_im = _RAND_2285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2286 = {1{`RANDOM}};
  _T_1312_re = _RAND_2286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2287 = {1{`RANDOM}};
  _T_1312_im = _RAND_2287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2288 = {1{`RANDOM}};
  _T_1313_re = _RAND_2288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2289 = {1{`RANDOM}};
  _T_1313_im = _RAND_2289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2290 = {1{`RANDOM}};
  _T_1314_re = _RAND_2290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2291 = {1{`RANDOM}};
  _T_1314_im = _RAND_2291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2292 = {1{`RANDOM}};
  _T_1315_re = _RAND_2292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2293 = {1{`RANDOM}};
  _T_1315_im = _RAND_2293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2294 = {1{`RANDOM}};
  _T_1316_re = _RAND_2294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2295 = {1{`RANDOM}};
  _T_1316_im = _RAND_2295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2296 = {1{`RANDOM}};
  _T_1317_re = _RAND_2296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2297 = {1{`RANDOM}};
  _T_1317_im = _RAND_2297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2298 = {1{`RANDOM}};
  _T_1318_re = _RAND_2298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2299 = {1{`RANDOM}};
  _T_1318_im = _RAND_2299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2300 = {1{`RANDOM}};
  _T_1319_re = _RAND_2300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2301 = {1{`RANDOM}};
  _T_1319_im = _RAND_2301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2302 = {1{`RANDOM}};
  _T_1320_re = _RAND_2302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2303 = {1{`RANDOM}};
  _T_1320_im = _RAND_2303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2304 = {1{`RANDOM}};
  _T_1321_re = _RAND_2304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2305 = {1{`RANDOM}};
  _T_1321_im = _RAND_2305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2306 = {1{`RANDOM}};
  _T_1327_re = _RAND_2306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2307 = {1{`RANDOM}};
  _T_1327_im = _RAND_2307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2308 = {1{`RANDOM}};
  _T_1328_re = _RAND_2308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2309 = {1{`RANDOM}};
  _T_1328_im = _RAND_2309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2310 = {1{`RANDOM}};
  _T_1329_re = _RAND_2310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2311 = {1{`RANDOM}};
  _T_1329_im = _RAND_2311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2312 = {1{`RANDOM}};
  _T_1330_re = _RAND_2312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2313 = {1{`RANDOM}};
  _T_1330_im = _RAND_2313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2314 = {1{`RANDOM}};
  _T_1331_re = _RAND_2314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2315 = {1{`RANDOM}};
  _T_1331_im = _RAND_2315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2316 = {1{`RANDOM}};
  _T_1332_re = _RAND_2316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2317 = {1{`RANDOM}};
  _T_1332_im = _RAND_2317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2318 = {1{`RANDOM}};
  _T_1333_re = _RAND_2318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2319 = {1{`RANDOM}};
  _T_1333_im = _RAND_2319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2320 = {1{`RANDOM}};
  _T_1334_re = _RAND_2320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2321 = {1{`RANDOM}};
  _T_1334_im = _RAND_2321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2322 = {1{`RANDOM}};
  _T_1335_re = _RAND_2322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2323 = {1{`RANDOM}};
  _T_1335_im = _RAND_2323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2324 = {1{`RANDOM}};
  _T_1336_re = _RAND_2324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2325 = {1{`RANDOM}};
  _T_1336_im = _RAND_2325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2326 = {1{`RANDOM}};
  _T_1337_re = _RAND_2326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2327 = {1{`RANDOM}};
  _T_1337_im = _RAND_2327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2328 = {1{`RANDOM}};
  _T_1338_re = _RAND_2328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2329 = {1{`RANDOM}};
  _T_1338_im = _RAND_2329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2330 = {1{`RANDOM}};
  _T_1339_re = _RAND_2330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2331 = {1{`RANDOM}};
  _T_1339_im = _RAND_2331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2332 = {1{`RANDOM}};
  _T_1340_re = _RAND_2332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2333 = {1{`RANDOM}};
  _T_1340_im = _RAND_2333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2334 = {1{`RANDOM}};
  _T_1341_re = _RAND_2334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2335 = {1{`RANDOM}};
  _T_1341_im = _RAND_2335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2336 = {1{`RANDOM}};
  _T_1342_re = _RAND_2336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2337 = {1{`RANDOM}};
  _T_1342_im = _RAND_2337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2338 = {1{`RANDOM}};
  _T_1343_re = _RAND_2338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2339 = {1{`RANDOM}};
  _T_1343_im = _RAND_2339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2340 = {1{`RANDOM}};
  _T_1344_re = _RAND_2340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2341 = {1{`RANDOM}};
  _T_1344_im = _RAND_2341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2342 = {1{`RANDOM}};
  _T_1345_re = _RAND_2342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2343 = {1{`RANDOM}};
  _T_1345_im = _RAND_2343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2344 = {1{`RANDOM}};
  _T_1346_re = _RAND_2344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2345 = {1{`RANDOM}};
  _T_1346_im = _RAND_2345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2346 = {1{`RANDOM}};
  _T_1347_re = _RAND_2346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2347 = {1{`RANDOM}};
  _T_1347_im = _RAND_2347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2348 = {1{`RANDOM}};
  _T_1348_re = _RAND_2348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2349 = {1{`RANDOM}};
  _T_1348_im = _RAND_2349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2350 = {1{`RANDOM}};
  _T_1349_re = _RAND_2350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2351 = {1{`RANDOM}};
  _T_1349_im = _RAND_2351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2352 = {1{`RANDOM}};
  _T_1350_re = _RAND_2352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2353 = {1{`RANDOM}};
  _T_1350_im = _RAND_2353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2354 = {1{`RANDOM}};
  _T_1351_re = _RAND_2354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2355 = {1{`RANDOM}};
  _T_1351_im = _RAND_2355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2356 = {1{`RANDOM}};
  _T_1352_re = _RAND_2356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2357 = {1{`RANDOM}};
  _T_1352_im = _RAND_2357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2358 = {1{`RANDOM}};
  _T_1353_re = _RAND_2358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2359 = {1{`RANDOM}};
  _T_1353_im = _RAND_2359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2360 = {1{`RANDOM}};
  _T_1354_re = _RAND_2360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2361 = {1{`RANDOM}};
  _T_1354_im = _RAND_2361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2362 = {1{`RANDOM}};
  _T_1355_re = _RAND_2362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2363 = {1{`RANDOM}};
  _T_1355_im = _RAND_2363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2364 = {1{`RANDOM}};
  _T_1356_re = _RAND_2364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2365 = {1{`RANDOM}};
  _T_1356_im = _RAND_2365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2366 = {1{`RANDOM}};
  _T_1357_re = _RAND_2366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2367 = {1{`RANDOM}};
  _T_1357_im = _RAND_2367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2368 = {1{`RANDOM}};
  _T_1358_re = _RAND_2368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2369 = {1{`RANDOM}};
  _T_1358_im = _RAND_2369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2370 = {1{`RANDOM}};
  _T_1359_re = _RAND_2370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2371 = {1{`RANDOM}};
  _T_1359_im = _RAND_2371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2372 = {1{`RANDOM}};
  _T_1360_re = _RAND_2372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2373 = {1{`RANDOM}};
  _T_1360_im = _RAND_2373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2374 = {1{`RANDOM}};
  _T_1361_re = _RAND_2374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2375 = {1{`RANDOM}};
  _T_1361_im = _RAND_2375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2376 = {1{`RANDOM}};
  _T_1362_re = _RAND_2376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2377 = {1{`RANDOM}};
  _T_1362_im = _RAND_2377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2378 = {1{`RANDOM}};
  _T_1363_re = _RAND_2378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2379 = {1{`RANDOM}};
  _T_1363_im = _RAND_2379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2380 = {1{`RANDOM}};
  _T_1364_re = _RAND_2380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2381 = {1{`RANDOM}};
  _T_1364_im = _RAND_2381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2382 = {1{`RANDOM}};
  _T_1365_re = _RAND_2382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2383 = {1{`RANDOM}};
  _T_1365_im = _RAND_2383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2384 = {1{`RANDOM}};
  _T_1366_re = _RAND_2384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2385 = {1{`RANDOM}};
  _T_1366_im = _RAND_2385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2386 = {1{`RANDOM}};
  _T_1367_re = _RAND_2386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2387 = {1{`RANDOM}};
  _T_1367_im = _RAND_2387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2388 = {1{`RANDOM}};
  _T_1368_re = _RAND_2388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2389 = {1{`RANDOM}};
  _T_1368_im = _RAND_2389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2390 = {1{`RANDOM}};
  _T_1369_re = _RAND_2390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2391 = {1{`RANDOM}};
  _T_1369_im = _RAND_2391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2392 = {1{`RANDOM}};
  _T_1370_re = _RAND_2392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2393 = {1{`RANDOM}};
  _T_1370_im = _RAND_2393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2394 = {1{`RANDOM}};
  _T_1371_re = _RAND_2394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2395 = {1{`RANDOM}};
  _T_1371_im = _RAND_2395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2396 = {1{`RANDOM}};
  _T_1372_re = _RAND_2396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2397 = {1{`RANDOM}};
  _T_1372_im = _RAND_2397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2398 = {1{`RANDOM}};
  _T_1373_re = _RAND_2398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2399 = {1{`RANDOM}};
  _T_1373_im = _RAND_2399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2400 = {1{`RANDOM}};
  _T_1374_re = _RAND_2400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2401 = {1{`RANDOM}};
  _T_1374_im = _RAND_2401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2402 = {1{`RANDOM}};
  _T_1375_re = _RAND_2402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2403 = {1{`RANDOM}};
  _T_1375_im = _RAND_2403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2404 = {1{`RANDOM}};
  _T_1376_re = _RAND_2404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2405 = {1{`RANDOM}};
  _T_1376_im = _RAND_2405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2406 = {1{`RANDOM}};
  _T_1377_re = _RAND_2406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2407 = {1{`RANDOM}};
  _T_1377_im = _RAND_2407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2408 = {1{`RANDOM}};
  _T_1378_re = _RAND_2408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2409 = {1{`RANDOM}};
  _T_1378_im = _RAND_2409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2410 = {1{`RANDOM}};
  _T_1379_re = _RAND_2410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2411 = {1{`RANDOM}};
  _T_1379_im = _RAND_2411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2412 = {1{`RANDOM}};
  _T_1380_re = _RAND_2412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2413 = {1{`RANDOM}};
  _T_1380_im = _RAND_2413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2414 = {1{`RANDOM}};
  _T_1381_re = _RAND_2414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2415 = {1{`RANDOM}};
  _T_1381_im = _RAND_2415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2416 = {1{`RANDOM}};
  _T_1382_re = _RAND_2416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2417 = {1{`RANDOM}};
  _T_1382_im = _RAND_2417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2418 = {1{`RANDOM}};
  _T_1383_re = _RAND_2418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2419 = {1{`RANDOM}};
  _T_1383_im = _RAND_2419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2420 = {1{`RANDOM}};
  _T_1384_re = _RAND_2420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2421 = {1{`RANDOM}};
  _T_1384_im = _RAND_2421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2422 = {1{`RANDOM}};
  _T_1385_re = _RAND_2422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2423 = {1{`RANDOM}};
  _T_1385_im = _RAND_2423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2424 = {1{`RANDOM}};
  _T_1386_re = _RAND_2424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2425 = {1{`RANDOM}};
  _T_1386_im = _RAND_2425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2426 = {1{`RANDOM}};
  _T_1387_re = _RAND_2426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2427 = {1{`RANDOM}};
  _T_1387_im = _RAND_2427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2428 = {1{`RANDOM}};
  _T_1388_re = _RAND_2428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2429 = {1{`RANDOM}};
  _T_1388_im = _RAND_2429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2430 = {1{`RANDOM}};
  _T_1389_re = _RAND_2430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2431 = {1{`RANDOM}};
  _T_1389_im = _RAND_2431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2432 = {1{`RANDOM}};
  _T_1390_re = _RAND_2432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2433 = {1{`RANDOM}};
  _T_1390_im = _RAND_2433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2434 = {1{`RANDOM}};
  _T_1391_re = _RAND_2434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2435 = {1{`RANDOM}};
  _T_1391_im = _RAND_2435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2436 = {1{`RANDOM}};
  _T_1392_re = _RAND_2436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2437 = {1{`RANDOM}};
  _T_1392_im = _RAND_2437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2438 = {1{`RANDOM}};
  _T_1393_re = _RAND_2438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2439 = {1{`RANDOM}};
  _T_1393_im = _RAND_2439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2440 = {1{`RANDOM}};
  _T_1394_re = _RAND_2440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2441 = {1{`RANDOM}};
  _T_1394_im = _RAND_2441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2442 = {1{`RANDOM}};
  _T_1395_re = _RAND_2442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2443 = {1{`RANDOM}};
  _T_1395_im = _RAND_2443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2444 = {1{`RANDOM}};
  _T_1396_re = _RAND_2444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2445 = {1{`RANDOM}};
  _T_1396_im = _RAND_2445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2446 = {1{`RANDOM}};
  _T_1397_re = _RAND_2446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2447 = {1{`RANDOM}};
  _T_1397_im = _RAND_2447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2448 = {1{`RANDOM}};
  _T_1398_re = _RAND_2448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2449 = {1{`RANDOM}};
  _T_1398_im = _RAND_2449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2450 = {1{`RANDOM}};
  _T_1399_re = _RAND_2450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2451 = {1{`RANDOM}};
  _T_1399_im = _RAND_2451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2452 = {1{`RANDOM}};
  _T_1400_re = _RAND_2452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2453 = {1{`RANDOM}};
  _T_1400_im = _RAND_2453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2454 = {1{`RANDOM}};
  _T_1401_re = _RAND_2454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2455 = {1{`RANDOM}};
  _T_1401_im = _RAND_2455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2456 = {1{`RANDOM}};
  _T_1402_re = _RAND_2456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2457 = {1{`RANDOM}};
  _T_1402_im = _RAND_2457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2458 = {1{`RANDOM}};
  _T_1403_re = _RAND_2458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2459 = {1{`RANDOM}};
  _T_1403_im = _RAND_2459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2460 = {1{`RANDOM}};
  _T_1404_re = _RAND_2460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2461 = {1{`RANDOM}};
  _T_1404_im = _RAND_2461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2462 = {1{`RANDOM}};
  _T_1405_re = _RAND_2462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2463 = {1{`RANDOM}};
  _T_1405_im = _RAND_2463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2464 = {1{`RANDOM}};
  _T_1406_re = _RAND_2464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2465 = {1{`RANDOM}};
  _T_1406_im = _RAND_2465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2466 = {1{`RANDOM}};
  _T_1407_re = _RAND_2466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2467 = {1{`RANDOM}};
  _T_1407_im = _RAND_2467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2468 = {1{`RANDOM}};
  _T_1408_re = _RAND_2468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2469 = {1{`RANDOM}};
  _T_1408_im = _RAND_2469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2470 = {1{`RANDOM}};
  _T_1409_re = _RAND_2470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2471 = {1{`RANDOM}};
  _T_1409_im = _RAND_2471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2472 = {1{`RANDOM}};
  _T_1410_re = _RAND_2472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2473 = {1{`RANDOM}};
  _T_1410_im = _RAND_2473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2474 = {1{`RANDOM}};
  _T_1411_re = _RAND_2474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2475 = {1{`RANDOM}};
  _T_1411_im = _RAND_2475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2476 = {1{`RANDOM}};
  _T_1412_re = _RAND_2476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2477 = {1{`RANDOM}};
  _T_1412_im = _RAND_2477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2478 = {1{`RANDOM}};
  _T_1413_re = _RAND_2478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2479 = {1{`RANDOM}};
  _T_1413_im = _RAND_2479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2480 = {1{`RANDOM}};
  _T_1414_re = _RAND_2480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2481 = {1{`RANDOM}};
  _T_1414_im = _RAND_2481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2482 = {1{`RANDOM}};
  _T_1415_re = _RAND_2482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2483 = {1{`RANDOM}};
  _T_1415_im = _RAND_2483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2484 = {1{`RANDOM}};
  _T_1416_re = _RAND_2484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2485 = {1{`RANDOM}};
  _T_1416_im = _RAND_2485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2486 = {1{`RANDOM}};
  _T_1417_re = _RAND_2486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2487 = {1{`RANDOM}};
  _T_1417_im = _RAND_2487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2488 = {1{`RANDOM}};
  _T_1418_re = _RAND_2488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2489 = {1{`RANDOM}};
  _T_1418_im = _RAND_2489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2490 = {1{`RANDOM}};
  _T_1419_re = _RAND_2490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2491 = {1{`RANDOM}};
  _T_1419_im = _RAND_2491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2492 = {1{`RANDOM}};
  _T_1420_re = _RAND_2492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2493 = {1{`RANDOM}};
  _T_1420_im = _RAND_2493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2494 = {1{`RANDOM}};
  _T_1421_re = _RAND_2494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2495 = {1{`RANDOM}};
  _T_1421_im = _RAND_2495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2496 = {1{`RANDOM}};
  _T_1422_re = _RAND_2496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2497 = {1{`RANDOM}};
  _T_1422_im = _RAND_2497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2498 = {1{`RANDOM}};
  _T_1423_re = _RAND_2498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2499 = {1{`RANDOM}};
  _T_1423_im = _RAND_2499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2500 = {1{`RANDOM}};
  _T_1424_re = _RAND_2500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2501 = {1{`RANDOM}};
  _T_1424_im = _RAND_2501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2502 = {1{`RANDOM}};
  _T_1425_re = _RAND_2502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2503 = {1{`RANDOM}};
  _T_1425_im = _RAND_2503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2504 = {1{`RANDOM}};
  _T_1426_re = _RAND_2504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2505 = {1{`RANDOM}};
  _T_1426_im = _RAND_2505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2506 = {1{`RANDOM}};
  _T_1427_re = _RAND_2506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2507 = {1{`RANDOM}};
  _T_1427_im = _RAND_2507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2508 = {1{`RANDOM}};
  _T_1428_re = _RAND_2508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2509 = {1{`RANDOM}};
  _T_1428_im = _RAND_2509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2510 = {1{`RANDOM}};
  _T_1429_re = _RAND_2510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2511 = {1{`RANDOM}};
  _T_1429_im = _RAND_2511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2512 = {1{`RANDOM}};
  _T_1430_re = _RAND_2512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2513 = {1{`RANDOM}};
  _T_1430_im = _RAND_2513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2514 = {1{`RANDOM}};
  _T_1431_re = _RAND_2514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2515 = {1{`RANDOM}};
  _T_1431_im = _RAND_2515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2516 = {1{`RANDOM}};
  _T_1432_re = _RAND_2516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2517 = {1{`RANDOM}};
  _T_1432_im = _RAND_2517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2518 = {1{`RANDOM}};
  _T_1433_re = _RAND_2518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2519 = {1{`RANDOM}};
  _T_1433_im = _RAND_2519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2520 = {1{`RANDOM}};
  _T_1434_re = _RAND_2520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2521 = {1{`RANDOM}};
  _T_1434_im = _RAND_2521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2522 = {1{`RANDOM}};
  _T_1435_re = _RAND_2522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2523 = {1{`RANDOM}};
  _T_1435_im = _RAND_2523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2524 = {1{`RANDOM}};
  _T_1436_re = _RAND_2524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2525 = {1{`RANDOM}};
  _T_1436_im = _RAND_2525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2526 = {1{`RANDOM}};
  _T_1437_re = _RAND_2526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2527 = {1{`RANDOM}};
  _T_1437_im = _RAND_2527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2528 = {1{`RANDOM}};
  _T_1438_re = _RAND_2528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2529 = {1{`RANDOM}};
  _T_1438_im = _RAND_2529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2530 = {1{`RANDOM}};
  _T_1439_re = _RAND_2530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2531 = {1{`RANDOM}};
  _T_1439_im = _RAND_2531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2532 = {1{`RANDOM}};
  _T_1440_re = _RAND_2532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2533 = {1{`RANDOM}};
  _T_1440_im = _RAND_2533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2534 = {1{`RANDOM}};
  _T_1441_re = _RAND_2534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2535 = {1{`RANDOM}};
  _T_1441_im = _RAND_2535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2536 = {1{`RANDOM}};
  _T_1442_re = _RAND_2536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2537 = {1{`RANDOM}};
  _T_1442_im = _RAND_2537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2538 = {1{`RANDOM}};
  _T_1443_re = _RAND_2538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2539 = {1{`RANDOM}};
  _T_1443_im = _RAND_2539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2540 = {1{`RANDOM}};
  _T_1444_re = _RAND_2540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2541 = {1{`RANDOM}};
  _T_1444_im = _RAND_2541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2542 = {1{`RANDOM}};
  _T_1445_re = _RAND_2542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2543 = {1{`RANDOM}};
  _T_1445_im = _RAND_2543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2544 = {1{`RANDOM}};
  _T_1446_re = _RAND_2544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2545 = {1{`RANDOM}};
  _T_1446_im = _RAND_2545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2546 = {1{`RANDOM}};
  _T_1447_re = _RAND_2546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2547 = {1{`RANDOM}};
  _T_1447_im = _RAND_2547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2548 = {1{`RANDOM}};
  _T_1448_re = _RAND_2548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2549 = {1{`RANDOM}};
  _T_1448_im = _RAND_2549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2550 = {1{`RANDOM}};
  _T_1449_re = _RAND_2550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2551 = {1{`RANDOM}};
  _T_1449_im = _RAND_2551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2552 = {1{`RANDOM}};
  _T_1450_re = _RAND_2552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2553 = {1{`RANDOM}};
  _T_1450_im = _RAND_2553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2554 = {1{`RANDOM}};
  _T_1451_re = _RAND_2554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2555 = {1{`RANDOM}};
  _T_1451_im = _RAND_2555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2556 = {1{`RANDOM}};
  _T_1452_re = _RAND_2556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2557 = {1{`RANDOM}};
  _T_1452_im = _RAND_2557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2558 = {1{`RANDOM}};
  _T_1453_re = _RAND_2558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2559 = {1{`RANDOM}};
  _T_1453_im = _RAND_2559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2560 = {1{`RANDOM}};
  _T_1454_re = _RAND_2560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2561 = {1{`RANDOM}};
  _T_1454_im = _RAND_2561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2562 = {1{`RANDOM}};
  _T_1457_re = _RAND_2562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2563 = {1{`RANDOM}};
  _T_1457_im = _RAND_2563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2564 = {1{`RANDOM}};
  _T_1458_re = _RAND_2564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2565 = {1{`RANDOM}};
  _T_1458_im = _RAND_2565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2566 = {1{`RANDOM}};
  _T_1459_re = _RAND_2566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2567 = {1{`RANDOM}};
  _T_1459_im = _RAND_2567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2568 = {1{`RANDOM}};
  _T_1460_re = _RAND_2568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2569 = {1{`RANDOM}};
  _T_1460_im = _RAND_2569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2570 = {1{`RANDOM}};
  _T_1461_re = _RAND_2570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2571 = {1{`RANDOM}};
  _T_1461_im = _RAND_2571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2572 = {1{`RANDOM}};
  _T_1462_re = _RAND_2572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2573 = {1{`RANDOM}};
  _T_1462_im = _RAND_2573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2574 = {1{`RANDOM}};
  _T_1463_re = _RAND_2574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2575 = {1{`RANDOM}};
  _T_1463_im = _RAND_2575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2576 = {1{`RANDOM}};
  _T_1464_re = _RAND_2576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2577 = {1{`RANDOM}};
  _T_1464_im = _RAND_2577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2578 = {1{`RANDOM}};
  _T_1465_re = _RAND_2578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2579 = {1{`RANDOM}};
  _T_1465_im = _RAND_2579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2580 = {1{`RANDOM}};
  _T_1466_re = _RAND_2580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2581 = {1{`RANDOM}};
  _T_1466_im = _RAND_2581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2582 = {1{`RANDOM}};
  _T_1467_re = _RAND_2582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2583 = {1{`RANDOM}};
  _T_1467_im = _RAND_2583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2584 = {1{`RANDOM}};
  _T_1468_re = _RAND_2584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2585 = {1{`RANDOM}};
  _T_1468_im = _RAND_2585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2586 = {1{`RANDOM}};
  _T_1469_re = _RAND_2586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2587 = {1{`RANDOM}};
  _T_1469_im = _RAND_2587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2588 = {1{`RANDOM}};
  _T_1470_re = _RAND_2588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2589 = {1{`RANDOM}};
  _T_1470_im = _RAND_2589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2590 = {1{`RANDOM}};
  _T_1471_re = _RAND_2590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2591 = {1{`RANDOM}};
  _T_1471_im = _RAND_2591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2592 = {1{`RANDOM}};
  _T_1472_re = _RAND_2592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2593 = {1{`RANDOM}};
  _T_1472_im = _RAND_2593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2594 = {1{`RANDOM}};
  _T_1473_re = _RAND_2594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2595 = {1{`RANDOM}};
  _T_1473_im = _RAND_2595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2596 = {1{`RANDOM}};
  _T_1474_re = _RAND_2596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2597 = {1{`RANDOM}};
  _T_1474_im = _RAND_2597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2598 = {1{`RANDOM}};
  _T_1475_re = _RAND_2598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2599 = {1{`RANDOM}};
  _T_1475_im = _RAND_2599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2600 = {1{`RANDOM}};
  _T_1476_re = _RAND_2600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2601 = {1{`RANDOM}};
  _T_1476_im = _RAND_2601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2602 = {1{`RANDOM}};
  _T_1477_re = _RAND_2602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2603 = {1{`RANDOM}};
  _T_1477_im = _RAND_2603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2604 = {1{`RANDOM}};
  _T_1478_re = _RAND_2604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2605 = {1{`RANDOM}};
  _T_1478_im = _RAND_2605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2606 = {1{`RANDOM}};
  _T_1479_re = _RAND_2606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2607 = {1{`RANDOM}};
  _T_1479_im = _RAND_2607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2608 = {1{`RANDOM}};
  _T_1480_re = _RAND_2608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2609 = {1{`RANDOM}};
  _T_1480_im = _RAND_2609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2610 = {1{`RANDOM}};
  _T_1481_re = _RAND_2610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2611 = {1{`RANDOM}};
  _T_1481_im = _RAND_2611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2612 = {1{`RANDOM}};
  _T_1482_re = _RAND_2612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2613 = {1{`RANDOM}};
  _T_1482_im = _RAND_2613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2614 = {1{`RANDOM}};
  _T_1483_re = _RAND_2614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2615 = {1{`RANDOM}};
  _T_1483_im = _RAND_2615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2616 = {1{`RANDOM}};
  _T_1484_re = _RAND_2616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2617 = {1{`RANDOM}};
  _T_1484_im = _RAND_2617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2618 = {1{`RANDOM}};
  _T_1485_re = _RAND_2618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2619 = {1{`RANDOM}};
  _T_1485_im = _RAND_2619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2620 = {1{`RANDOM}};
  _T_1486_re = _RAND_2620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2621 = {1{`RANDOM}};
  _T_1486_im = _RAND_2621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2622 = {1{`RANDOM}};
  _T_1487_re = _RAND_2622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2623 = {1{`RANDOM}};
  _T_1487_im = _RAND_2623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2624 = {1{`RANDOM}};
  _T_1488_re = _RAND_2624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2625 = {1{`RANDOM}};
  _T_1488_im = _RAND_2625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2626 = {1{`RANDOM}};
  _T_1489_re = _RAND_2626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2627 = {1{`RANDOM}};
  _T_1489_im = _RAND_2627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2628 = {1{`RANDOM}};
  _T_1490_re = _RAND_2628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2629 = {1{`RANDOM}};
  _T_1490_im = _RAND_2629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2630 = {1{`RANDOM}};
  _T_1491_re = _RAND_2630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2631 = {1{`RANDOM}};
  _T_1491_im = _RAND_2631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2632 = {1{`RANDOM}};
  _T_1492_re = _RAND_2632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2633 = {1{`RANDOM}};
  _T_1492_im = _RAND_2633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2634 = {1{`RANDOM}};
  _T_1493_re = _RAND_2634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2635 = {1{`RANDOM}};
  _T_1493_im = _RAND_2635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2636 = {1{`RANDOM}};
  _T_1494_re = _RAND_2636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2637 = {1{`RANDOM}};
  _T_1494_im = _RAND_2637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2638 = {1{`RANDOM}};
  _T_1495_re = _RAND_2638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2639 = {1{`RANDOM}};
  _T_1495_im = _RAND_2639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2640 = {1{`RANDOM}};
  _T_1496_re = _RAND_2640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2641 = {1{`RANDOM}};
  _T_1496_im = _RAND_2641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2642 = {1{`RANDOM}};
  _T_1497_re = _RAND_2642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2643 = {1{`RANDOM}};
  _T_1497_im = _RAND_2643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2644 = {1{`RANDOM}};
  _T_1498_re = _RAND_2644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2645 = {1{`RANDOM}};
  _T_1498_im = _RAND_2645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2646 = {1{`RANDOM}};
  _T_1499_re = _RAND_2646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2647 = {1{`RANDOM}};
  _T_1499_im = _RAND_2647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2648 = {1{`RANDOM}};
  _T_1500_re = _RAND_2648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2649 = {1{`RANDOM}};
  _T_1500_im = _RAND_2649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2650 = {1{`RANDOM}};
  _T_1501_re = _RAND_2650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2651 = {1{`RANDOM}};
  _T_1501_im = _RAND_2651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2652 = {1{`RANDOM}};
  _T_1502_re = _RAND_2652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2653 = {1{`RANDOM}};
  _T_1502_im = _RAND_2653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2654 = {1{`RANDOM}};
  _T_1503_re = _RAND_2654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2655 = {1{`RANDOM}};
  _T_1503_im = _RAND_2655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2656 = {1{`RANDOM}};
  _T_1504_re = _RAND_2656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2657 = {1{`RANDOM}};
  _T_1504_im = _RAND_2657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2658 = {1{`RANDOM}};
  _T_1505_re = _RAND_2658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2659 = {1{`RANDOM}};
  _T_1505_im = _RAND_2659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2660 = {1{`RANDOM}};
  _T_1506_re = _RAND_2660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2661 = {1{`RANDOM}};
  _T_1506_im = _RAND_2661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2662 = {1{`RANDOM}};
  _T_1507_re = _RAND_2662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2663 = {1{`RANDOM}};
  _T_1507_im = _RAND_2663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2664 = {1{`RANDOM}};
  _T_1508_re = _RAND_2664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2665 = {1{`RANDOM}};
  _T_1508_im = _RAND_2665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2666 = {1{`RANDOM}};
  _T_1509_re = _RAND_2666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2667 = {1{`RANDOM}};
  _T_1509_im = _RAND_2667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2668 = {1{`RANDOM}};
  _T_1510_re = _RAND_2668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2669 = {1{`RANDOM}};
  _T_1510_im = _RAND_2669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2670 = {1{`RANDOM}};
  _T_1511_re = _RAND_2670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2671 = {1{`RANDOM}};
  _T_1511_im = _RAND_2671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2672 = {1{`RANDOM}};
  _T_1512_re = _RAND_2672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2673 = {1{`RANDOM}};
  _T_1512_im = _RAND_2673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2674 = {1{`RANDOM}};
  _T_1513_re = _RAND_2674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2675 = {1{`RANDOM}};
  _T_1513_im = _RAND_2675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2676 = {1{`RANDOM}};
  _T_1514_re = _RAND_2676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2677 = {1{`RANDOM}};
  _T_1514_im = _RAND_2677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2678 = {1{`RANDOM}};
  _T_1515_re = _RAND_2678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2679 = {1{`RANDOM}};
  _T_1515_im = _RAND_2679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2680 = {1{`RANDOM}};
  _T_1516_re = _RAND_2680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2681 = {1{`RANDOM}};
  _T_1516_im = _RAND_2681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2682 = {1{`RANDOM}};
  _T_1517_re = _RAND_2682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2683 = {1{`RANDOM}};
  _T_1517_im = _RAND_2683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2684 = {1{`RANDOM}};
  _T_1518_re = _RAND_2684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2685 = {1{`RANDOM}};
  _T_1518_im = _RAND_2685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2686 = {1{`RANDOM}};
  _T_1519_re = _RAND_2686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2687 = {1{`RANDOM}};
  _T_1519_im = _RAND_2687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2688 = {1{`RANDOM}};
  _T_1520_re = _RAND_2688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2689 = {1{`RANDOM}};
  _T_1520_im = _RAND_2689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2690 = {1{`RANDOM}};
  _T_1526_re = _RAND_2690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2691 = {1{`RANDOM}};
  _T_1526_im = _RAND_2691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2692 = {1{`RANDOM}};
  _T_1527_re = _RAND_2692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2693 = {1{`RANDOM}};
  _T_1527_im = _RAND_2693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2694 = {1{`RANDOM}};
  _T_1528_re = _RAND_2694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2695 = {1{`RANDOM}};
  _T_1528_im = _RAND_2695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2696 = {1{`RANDOM}};
  _T_1529_re = _RAND_2696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2697 = {1{`RANDOM}};
  _T_1529_im = _RAND_2697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2698 = {1{`RANDOM}};
  _T_1530_re = _RAND_2698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2699 = {1{`RANDOM}};
  _T_1530_im = _RAND_2699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2700 = {1{`RANDOM}};
  _T_1531_re = _RAND_2700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2701 = {1{`RANDOM}};
  _T_1531_im = _RAND_2701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2702 = {1{`RANDOM}};
  _T_1532_re = _RAND_2702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2703 = {1{`RANDOM}};
  _T_1532_im = _RAND_2703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2704 = {1{`RANDOM}};
  _T_1533_re = _RAND_2704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2705 = {1{`RANDOM}};
  _T_1533_im = _RAND_2705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2706 = {1{`RANDOM}};
  _T_1534_re = _RAND_2706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2707 = {1{`RANDOM}};
  _T_1534_im = _RAND_2707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2708 = {1{`RANDOM}};
  _T_1535_re = _RAND_2708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2709 = {1{`RANDOM}};
  _T_1535_im = _RAND_2709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2710 = {1{`RANDOM}};
  _T_1536_re = _RAND_2710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2711 = {1{`RANDOM}};
  _T_1536_im = _RAND_2711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2712 = {1{`RANDOM}};
  _T_1537_re = _RAND_2712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2713 = {1{`RANDOM}};
  _T_1537_im = _RAND_2713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2714 = {1{`RANDOM}};
  _T_1538_re = _RAND_2714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2715 = {1{`RANDOM}};
  _T_1538_im = _RAND_2715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2716 = {1{`RANDOM}};
  _T_1539_re = _RAND_2716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2717 = {1{`RANDOM}};
  _T_1539_im = _RAND_2717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2718 = {1{`RANDOM}};
  _T_1540_re = _RAND_2718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2719 = {1{`RANDOM}};
  _T_1540_im = _RAND_2719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2720 = {1{`RANDOM}};
  _T_1541_re = _RAND_2720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2721 = {1{`RANDOM}};
  _T_1541_im = _RAND_2721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2722 = {1{`RANDOM}};
  _T_1542_re = _RAND_2722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2723 = {1{`RANDOM}};
  _T_1542_im = _RAND_2723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2724 = {1{`RANDOM}};
  _T_1543_re = _RAND_2724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2725 = {1{`RANDOM}};
  _T_1543_im = _RAND_2725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2726 = {1{`RANDOM}};
  _T_1544_re = _RAND_2726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2727 = {1{`RANDOM}};
  _T_1544_im = _RAND_2727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2728 = {1{`RANDOM}};
  _T_1545_re = _RAND_2728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2729 = {1{`RANDOM}};
  _T_1545_im = _RAND_2729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2730 = {1{`RANDOM}};
  _T_1546_re = _RAND_2730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2731 = {1{`RANDOM}};
  _T_1546_im = _RAND_2731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2732 = {1{`RANDOM}};
  _T_1547_re = _RAND_2732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2733 = {1{`RANDOM}};
  _T_1547_im = _RAND_2733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2734 = {1{`RANDOM}};
  _T_1548_re = _RAND_2734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2735 = {1{`RANDOM}};
  _T_1548_im = _RAND_2735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2736 = {1{`RANDOM}};
  _T_1549_re = _RAND_2736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2737 = {1{`RANDOM}};
  _T_1549_im = _RAND_2737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2738 = {1{`RANDOM}};
  _T_1550_re = _RAND_2738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2739 = {1{`RANDOM}};
  _T_1550_im = _RAND_2739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2740 = {1{`RANDOM}};
  _T_1551_re = _RAND_2740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2741 = {1{`RANDOM}};
  _T_1551_im = _RAND_2741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2742 = {1{`RANDOM}};
  _T_1552_re = _RAND_2742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2743 = {1{`RANDOM}};
  _T_1552_im = _RAND_2743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2744 = {1{`RANDOM}};
  _T_1553_re = _RAND_2744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2745 = {1{`RANDOM}};
  _T_1553_im = _RAND_2745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2746 = {1{`RANDOM}};
  _T_1554_re = _RAND_2746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2747 = {1{`RANDOM}};
  _T_1554_im = _RAND_2747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2748 = {1{`RANDOM}};
  _T_1555_re = _RAND_2748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2749 = {1{`RANDOM}};
  _T_1555_im = _RAND_2749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2750 = {1{`RANDOM}};
  _T_1556_re = _RAND_2750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2751 = {1{`RANDOM}};
  _T_1556_im = _RAND_2751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2752 = {1{`RANDOM}};
  _T_1557_re = _RAND_2752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2753 = {1{`RANDOM}};
  _T_1557_im = _RAND_2753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2754 = {1{`RANDOM}};
  _T_1558_re = _RAND_2754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2755 = {1{`RANDOM}};
  _T_1558_im = _RAND_2755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2756 = {1{`RANDOM}};
  _T_1559_re = _RAND_2756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2757 = {1{`RANDOM}};
  _T_1559_im = _RAND_2757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2758 = {1{`RANDOM}};
  _T_1560_re = _RAND_2758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2759 = {1{`RANDOM}};
  _T_1560_im = _RAND_2759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2760 = {1{`RANDOM}};
  _T_1561_re = _RAND_2760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2761 = {1{`RANDOM}};
  _T_1561_im = _RAND_2761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2762 = {1{`RANDOM}};
  _T_1562_re = _RAND_2762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2763 = {1{`RANDOM}};
  _T_1562_im = _RAND_2763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2764 = {1{`RANDOM}};
  _T_1563_re = _RAND_2764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2765 = {1{`RANDOM}};
  _T_1563_im = _RAND_2765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2766 = {1{`RANDOM}};
  _T_1564_re = _RAND_2766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2767 = {1{`RANDOM}};
  _T_1564_im = _RAND_2767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2768 = {1{`RANDOM}};
  _T_1565_re = _RAND_2768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2769 = {1{`RANDOM}};
  _T_1565_im = _RAND_2769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2770 = {1{`RANDOM}};
  _T_1566_re = _RAND_2770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2771 = {1{`RANDOM}};
  _T_1566_im = _RAND_2771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2772 = {1{`RANDOM}};
  _T_1567_re = _RAND_2772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2773 = {1{`RANDOM}};
  _T_1567_im = _RAND_2773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2774 = {1{`RANDOM}};
  _T_1568_re = _RAND_2774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2775 = {1{`RANDOM}};
  _T_1568_im = _RAND_2775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2776 = {1{`RANDOM}};
  _T_1569_re = _RAND_2776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2777 = {1{`RANDOM}};
  _T_1569_im = _RAND_2777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2778 = {1{`RANDOM}};
  _T_1570_re = _RAND_2778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2779 = {1{`RANDOM}};
  _T_1570_im = _RAND_2779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2780 = {1{`RANDOM}};
  _T_1571_re = _RAND_2780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2781 = {1{`RANDOM}};
  _T_1571_im = _RAND_2781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2782 = {1{`RANDOM}};
  _T_1572_re = _RAND_2782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2783 = {1{`RANDOM}};
  _T_1572_im = _RAND_2783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2784 = {1{`RANDOM}};
  _T_1573_re = _RAND_2784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2785 = {1{`RANDOM}};
  _T_1573_im = _RAND_2785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2786 = {1{`RANDOM}};
  _T_1574_re = _RAND_2786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2787 = {1{`RANDOM}};
  _T_1574_im = _RAND_2787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2788 = {1{`RANDOM}};
  _T_1575_re = _RAND_2788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2789 = {1{`RANDOM}};
  _T_1575_im = _RAND_2789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2790 = {1{`RANDOM}};
  _T_1576_re = _RAND_2790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2791 = {1{`RANDOM}};
  _T_1576_im = _RAND_2791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2792 = {1{`RANDOM}};
  _T_1577_re = _RAND_2792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2793 = {1{`RANDOM}};
  _T_1577_im = _RAND_2793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2794 = {1{`RANDOM}};
  _T_1578_re = _RAND_2794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2795 = {1{`RANDOM}};
  _T_1578_im = _RAND_2795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2796 = {1{`RANDOM}};
  _T_1579_re = _RAND_2796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2797 = {1{`RANDOM}};
  _T_1579_im = _RAND_2797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2798 = {1{`RANDOM}};
  _T_1580_re = _RAND_2798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2799 = {1{`RANDOM}};
  _T_1580_im = _RAND_2799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2800 = {1{`RANDOM}};
  _T_1581_re = _RAND_2800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2801 = {1{`RANDOM}};
  _T_1581_im = _RAND_2801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2802 = {1{`RANDOM}};
  _T_1582_re = _RAND_2802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2803 = {1{`RANDOM}};
  _T_1582_im = _RAND_2803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2804 = {1{`RANDOM}};
  _T_1583_re = _RAND_2804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2805 = {1{`RANDOM}};
  _T_1583_im = _RAND_2805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2806 = {1{`RANDOM}};
  _T_1584_re = _RAND_2806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2807 = {1{`RANDOM}};
  _T_1584_im = _RAND_2807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2808 = {1{`RANDOM}};
  _T_1585_re = _RAND_2808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2809 = {1{`RANDOM}};
  _T_1585_im = _RAND_2809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2810 = {1{`RANDOM}};
  _T_1586_re = _RAND_2810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2811 = {1{`RANDOM}};
  _T_1586_im = _RAND_2811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2812 = {1{`RANDOM}};
  _T_1587_re = _RAND_2812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2813 = {1{`RANDOM}};
  _T_1587_im = _RAND_2813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2814 = {1{`RANDOM}};
  _T_1588_re = _RAND_2814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2815 = {1{`RANDOM}};
  _T_1588_im = _RAND_2815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2816 = {1{`RANDOM}};
  _T_1589_re = _RAND_2816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2817 = {1{`RANDOM}};
  _T_1589_im = _RAND_2817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2818 = {1{`RANDOM}};
  _T_1592_re = _RAND_2818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2819 = {1{`RANDOM}};
  _T_1592_im = _RAND_2819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2820 = {1{`RANDOM}};
  _T_1593_re = _RAND_2820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2821 = {1{`RANDOM}};
  _T_1593_im = _RAND_2821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2822 = {1{`RANDOM}};
  _T_1594_re = _RAND_2822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2823 = {1{`RANDOM}};
  _T_1594_im = _RAND_2823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2824 = {1{`RANDOM}};
  _T_1595_re = _RAND_2824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2825 = {1{`RANDOM}};
  _T_1595_im = _RAND_2825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2826 = {1{`RANDOM}};
  _T_1596_re = _RAND_2826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2827 = {1{`RANDOM}};
  _T_1596_im = _RAND_2827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2828 = {1{`RANDOM}};
  _T_1597_re = _RAND_2828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2829 = {1{`RANDOM}};
  _T_1597_im = _RAND_2829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2830 = {1{`RANDOM}};
  _T_1598_re = _RAND_2830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2831 = {1{`RANDOM}};
  _T_1598_im = _RAND_2831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2832 = {1{`RANDOM}};
  _T_1599_re = _RAND_2832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2833 = {1{`RANDOM}};
  _T_1599_im = _RAND_2833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2834 = {1{`RANDOM}};
  _T_1600_re = _RAND_2834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2835 = {1{`RANDOM}};
  _T_1600_im = _RAND_2835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2836 = {1{`RANDOM}};
  _T_1601_re = _RAND_2836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2837 = {1{`RANDOM}};
  _T_1601_im = _RAND_2837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2838 = {1{`RANDOM}};
  _T_1602_re = _RAND_2838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2839 = {1{`RANDOM}};
  _T_1602_im = _RAND_2839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2840 = {1{`RANDOM}};
  _T_1603_re = _RAND_2840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2841 = {1{`RANDOM}};
  _T_1603_im = _RAND_2841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2842 = {1{`RANDOM}};
  _T_1604_re = _RAND_2842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2843 = {1{`RANDOM}};
  _T_1604_im = _RAND_2843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2844 = {1{`RANDOM}};
  _T_1605_re = _RAND_2844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2845 = {1{`RANDOM}};
  _T_1605_im = _RAND_2845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2846 = {1{`RANDOM}};
  _T_1606_re = _RAND_2846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2847 = {1{`RANDOM}};
  _T_1606_im = _RAND_2847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2848 = {1{`RANDOM}};
  _T_1607_re = _RAND_2848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2849 = {1{`RANDOM}};
  _T_1607_im = _RAND_2849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2850 = {1{`RANDOM}};
  _T_1608_re = _RAND_2850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2851 = {1{`RANDOM}};
  _T_1608_im = _RAND_2851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2852 = {1{`RANDOM}};
  _T_1609_re = _RAND_2852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2853 = {1{`RANDOM}};
  _T_1609_im = _RAND_2853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2854 = {1{`RANDOM}};
  _T_1610_re = _RAND_2854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2855 = {1{`RANDOM}};
  _T_1610_im = _RAND_2855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2856 = {1{`RANDOM}};
  _T_1611_re = _RAND_2856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2857 = {1{`RANDOM}};
  _T_1611_im = _RAND_2857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2858 = {1{`RANDOM}};
  _T_1612_re = _RAND_2858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2859 = {1{`RANDOM}};
  _T_1612_im = _RAND_2859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2860 = {1{`RANDOM}};
  _T_1613_re = _RAND_2860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2861 = {1{`RANDOM}};
  _T_1613_im = _RAND_2861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2862 = {1{`RANDOM}};
  _T_1614_re = _RAND_2862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2863 = {1{`RANDOM}};
  _T_1614_im = _RAND_2863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2864 = {1{`RANDOM}};
  _T_1615_re = _RAND_2864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2865 = {1{`RANDOM}};
  _T_1615_im = _RAND_2865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2866 = {1{`RANDOM}};
  _T_1616_re = _RAND_2866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2867 = {1{`RANDOM}};
  _T_1616_im = _RAND_2867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2868 = {1{`RANDOM}};
  _T_1617_re = _RAND_2868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2869 = {1{`RANDOM}};
  _T_1617_im = _RAND_2869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2870 = {1{`RANDOM}};
  _T_1618_re = _RAND_2870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2871 = {1{`RANDOM}};
  _T_1618_im = _RAND_2871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2872 = {1{`RANDOM}};
  _T_1619_re = _RAND_2872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2873 = {1{`RANDOM}};
  _T_1619_im = _RAND_2873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2874 = {1{`RANDOM}};
  _T_1620_re = _RAND_2874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2875 = {1{`RANDOM}};
  _T_1620_im = _RAND_2875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2876 = {1{`RANDOM}};
  _T_1621_re = _RAND_2876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2877 = {1{`RANDOM}};
  _T_1621_im = _RAND_2877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2878 = {1{`RANDOM}};
  _T_1622_re = _RAND_2878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2879 = {1{`RANDOM}};
  _T_1622_im = _RAND_2879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2880 = {1{`RANDOM}};
  _T_1623_re = _RAND_2880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2881 = {1{`RANDOM}};
  _T_1623_im = _RAND_2881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2882 = {1{`RANDOM}};
  _T_1629_re = _RAND_2882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2883 = {1{`RANDOM}};
  _T_1629_im = _RAND_2883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2884 = {1{`RANDOM}};
  _T_1630_re = _RAND_2884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2885 = {1{`RANDOM}};
  _T_1630_im = _RAND_2885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2886 = {1{`RANDOM}};
  _T_1631_re = _RAND_2886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2887 = {1{`RANDOM}};
  _T_1631_im = _RAND_2887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2888 = {1{`RANDOM}};
  _T_1632_re = _RAND_2888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2889 = {1{`RANDOM}};
  _T_1632_im = _RAND_2889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2890 = {1{`RANDOM}};
  _T_1633_re = _RAND_2890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2891 = {1{`RANDOM}};
  _T_1633_im = _RAND_2891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2892 = {1{`RANDOM}};
  _T_1634_re = _RAND_2892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2893 = {1{`RANDOM}};
  _T_1634_im = _RAND_2893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2894 = {1{`RANDOM}};
  _T_1635_re = _RAND_2894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2895 = {1{`RANDOM}};
  _T_1635_im = _RAND_2895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2896 = {1{`RANDOM}};
  _T_1636_re = _RAND_2896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2897 = {1{`RANDOM}};
  _T_1636_im = _RAND_2897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2898 = {1{`RANDOM}};
  _T_1637_re = _RAND_2898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2899 = {1{`RANDOM}};
  _T_1637_im = _RAND_2899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2900 = {1{`RANDOM}};
  _T_1638_re = _RAND_2900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2901 = {1{`RANDOM}};
  _T_1638_im = _RAND_2901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2902 = {1{`RANDOM}};
  _T_1639_re = _RAND_2902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2903 = {1{`RANDOM}};
  _T_1639_im = _RAND_2903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2904 = {1{`RANDOM}};
  _T_1640_re = _RAND_2904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2905 = {1{`RANDOM}};
  _T_1640_im = _RAND_2905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2906 = {1{`RANDOM}};
  _T_1641_re = _RAND_2906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2907 = {1{`RANDOM}};
  _T_1641_im = _RAND_2907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2908 = {1{`RANDOM}};
  _T_1642_re = _RAND_2908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2909 = {1{`RANDOM}};
  _T_1642_im = _RAND_2909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2910 = {1{`RANDOM}};
  _T_1643_re = _RAND_2910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2911 = {1{`RANDOM}};
  _T_1643_im = _RAND_2911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2912 = {1{`RANDOM}};
  _T_1644_re = _RAND_2912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2913 = {1{`RANDOM}};
  _T_1644_im = _RAND_2913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2914 = {1{`RANDOM}};
  _T_1645_re = _RAND_2914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2915 = {1{`RANDOM}};
  _T_1645_im = _RAND_2915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2916 = {1{`RANDOM}};
  _T_1646_re = _RAND_2916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2917 = {1{`RANDOM}};
  _T_1646_im = _RAND_2917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2918 = {1{`RANDOM}};
  _T_1647_re = _RAND_2918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2919 = {1{`RANDOM}};
  _T_1647_im = _RAND_2919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2920 = {1{`RANDOM}};
  _T_1648_re = _RAND_2920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2921 = {1{`RANDOM}};
  _T_1648_im = _RAND_2921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2922 = {1{`RANDOM}};
  _T_1649_re = _RAND_2922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2923 = {1{`RANDOM}};
  _T_1649_im = _RAND_2923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2924 = {1{`RANDOM}};
  _T_1650_re = _RAND_2924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2925 = {1{`RANDOM}};
  _T_1650_im = _RAND_2925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2926 = {1{`RANDOM}};
  _T_1651_re = _RAND_2926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2927 = {1{`RANDOM}};
  _T_1651_im = _RAND_2927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2928 = {1{`RANDOM}};
  _T_1652_re = _RAND_2928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2929 = {1{`RANDOM}};
  _T_1652_im = _RAND_2929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2930 = {1{`RANDOM}};
  _T_1653_re = _RAND_2930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2931 = {1{`RANDOM}};
  _T_1653_im = _RAND_2931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2932 = {1{`RANDOM}};
  _T_1654_re = _RAND_2932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2933 = {1{`RANDOM}};
  _T_1654_im = _RAND_2933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2934 = {1{`RANDOM}};
  _T_1655_re = _RAND_2934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2935 = {1{`RANDOM}};
  _T_1655_im = _RAND_2935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2936 = {1{`RANDOM}};
  _T_1656_re = _RAND_2936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2937 = {1{`RANDOM}};
  _T_1656_im = _RAND_2937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2938 = {1{`RANDOM}};
  _T_1657_re = _RAND_2938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2939 = {1{`RANDOM}};
  _T_1657_im = _RAND_2939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2940 = {1{`RANDOM}};
  _T_1658_re = _RAND_2940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2941 = {1{`RANDOM}};
  _T_1658_im = _RAND_2941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2942 = {1{`RANDOM}};
  _T_1659_re = _RAND_2942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2943 = {1{`RANDOM}};
  _T_1659_im = _RAND_2943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2944 = {1{`RANDOM}};
  _T_1660_re = _RAND_2944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2945 = {1{`RANDOM}};
  _T_1660_im = _RAND_2945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2946 = {1{`RANDOM}};
  _T_1663_re = _RAND_2946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2947 = {1{`RANDOM}};
  _T_1663_im = _RAND_2947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2948 = {1{`RANDOM}};
  _T_1664_re = _RAND_2948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2949 = {1{`RANDOM}};
  _T_1664_im = _RAND_2949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2950 = {1{`RANDOM}};
  _T_1665_re = _RAND_2950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2951 = {1{`RANDOM}};
  _T_1665_im = _RAND_2951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2952 = {1{`RANDOM}};
  _T_1666_re = _RAND_2952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2953 = {1{`RANDOM}};
  _T_1666_im = _RAND_2953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2954 = {1{`RANDOM}};
  _T_1667_re = _RAND_2954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2955 = {1{`RANDOM}};
  _T_1667_im = _RAND_2955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2956 = {1{`RANDOM}};
  _T_1668_re = _RAND_2956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2957 = {1{`RANDOM}};
  _T_1668_im = _RAND_2957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2958 = {1{`RANDOM}};
  _T_1669_re = _RAND_2958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2959 = {1{`RANDOM}};
  _T_1669_im = _RAND_2959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2960 = {1{`RANDOM}};
  _T_1670_re = _RAND_2960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2961 = {1{`RANDOM}};
  _T_1670_im = _RAND_2961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2962 = {1{`RANDOM}};
  _T_1671_re = _RAND_2962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2963 = {1{`RANDOM}};
  _T_1671_im = _RAND_2963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2964 = {1{`RANDOM}};
  _T_1672_re = _RAND_2964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2965 = {1{`RANDOM}};
  _T_1672_im = _RAND_2965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2966 = {1{`RANDOM}};
  _T_1673_re = _RAND_2966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2967 = {1{`RANDOM}};
  _T_1673_im = _RAND_2967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2968 = {1{`RANDOM}};
  _T_1674_re = _RAND_2968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2969 = {1{`RANDOM}};
  _T_1674_im = _RAND_2969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2970 = {1{`RANDOM}};
  _T_1675_re = _RAND_2970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2971 = {1{`RANDOM}};
  _T_1675_im = _RAND_2971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2972 = {1{`RANDOM}};
  _T_1676_re = _RAND_2972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2973 = {1{`RANDOM}};
  _T_1676_im = _RAND_2973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2974 = {1{`RANDOM}};
  _T_1677_re = _RAND_2974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2975 = {1{`RANDOM}};
  _T_1677_im = _RAND_2975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2976 = {1{`RANDOM}};
  _T_1678_re = _RAND_2976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2977 = {1{`RANDOM}};
  _T_1678_im = _RAND_2977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2978 = {1{`RANDOM}};
  _T_1684_re = _RAND_2978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2979 = {1{`RANDOM}};
  _T_1684_im = _RAND_2979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2980 = {1{`RANDOM}};
  _T_1685_re = _RAND_2980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2981 = {1{`RANDOM}};
  _T_1685_im = _RAND_2981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2982 = {1{`RANDOM}};
  _T_1686_re = _RAND_2982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2983 = {1{`RANDOM}};
  _T_1686_im = _RAND_2983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2984 = {1{`RANDOM}};
  _T_1687_re = _RAND_2984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2985 = {1{`RANDOM}};
  _T_1687_im = _RAND_2985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2986 = {1{`RANDOM}};
  _T_1688_re = _RAND_2986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2987 = {1{`RANDOM}};
  _T_1688_im = _RAND_2987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2988 = {1{`RANDOM}};
  _T_1689_re = _RAND_2988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2989 = {1{`RANDOM}};
  _T_1689_im = _RAND_2989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2990 = {1{`RANDOM}};
  _T_1690_re = _RAND_2990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2991 = {1{`RANDOM}};
  _T_1690_im = _RAND_2991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2992 = {1{`RANDOM}};
  _T_1691_re = _RAND_2992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2993 = {1{`RANDOM}};
  _T_1691_im = _RAND_2993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2994 = {1{`RANDOM}};
  _T_1692_re = _RAND_2994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2995 = {1{`RANDOM}};
  _T_1692_im = _RAND_2995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2996 = {1{`RANDOM}};
  _T_1693_re = _RAND_2996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2997 = {1{`RANDOM}};
  _T_1693_im = _RAND_2997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2998 = {1{`RANDOM}};
  _T_1694_re = _RAND_2998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2999 = {1{`RANDOM}};
  _T_1694_im = _RAND_2999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3000 = {1{`RANDOM}};
  _T_1695_re = _RAND_3000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3001 = {1{`RANDOM}};
  _T_1695_im = _RAND_3001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3002 = {1{`RANDOM}};
  _T_1696_re = _RAND_3002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3003 = {1{`RANDOM}};
  _T_1696_im = _RAND_3003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3004 = {1{`RANDOM}};
  _T_1697_re = _RAND_3004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3005 = {1{`RANDOM}};
  _T_1697_im = _RAND_3005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3006 = {1{`RANDOM}};
  _T_1698_re = _RAND_3006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3007 = {1{`RANDOM}};
  _T_1698_im = _RAND_3007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3008 = {1{`RANDOM}};
  _T_1699_re = _RAND_3008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3009 = {1{`RANDOM}};
  _T_1699_im = _RAND_3009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3010 = {1{`RANDOM}};
  _T_1702_re = _RAND_3010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3011 = {1{`RANDOM}};
  _T_1702_im = _RAND_3011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3012 = {1{`RANDOM}};
  _T_1703_re = _RAND_3012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3013 = {1{`RANDOM}};
  _T_1703_im = _RAND_3013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3014 = {1{`RANDOM}};
  _T_1704_re = _RAND_3014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3015 = {1{`RANDOM}};
  _T_1704_im = _RAND_3015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3016 = {1{`RANDOM}};
  _T_1705_re = _RAND_3016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3017 = {1{`RANDOM}};
  _T_1705_im = _RAND_3017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3018 = {1{`RANDOM}};
  _T_1706_re = _RAND_3018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3019 = {1{`RANDOM}};
  _T_1706_im = _RAND_3019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3020 = {1{`RANDOM}};
  _T_1707_re = _RAND_3020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3021 = {1{`RANDOM}};
  _T_1707_im = _RAND_3021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3022 = {1{`RANDOM}};
  _T_1708_re = _RAND_3022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3023 = {1{`RANDOM}};
  _T_1708_im = _RAND_3023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3024 = {1{`RANDOM}};
  _T_1709_re = _RAND_3024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3025 = {1{`RANDOM}};
  _T_1709_im = _RAND_3025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3026 = {1{`RANDOM}};
  _T_1715_re = _RAND_3026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3027 = {1{`RANDOM}};
  _T_1715_im = _RAND_3027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3028 = {1{`RANDOM}};
  _T_1716_re = _RAND_3028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3029 = {1{`RANDOM}};
  _T_1716_im = _RAND_3029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3030 = {1{`RANDOM}};
  _T_1717_re = _RAND_3030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3031 = {1{`RANDOM}};
  _T_1717_im = _RAND_3031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3032 = {1{`RANDOM}};
  _T_1718_re = _RAND_3032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3033 = {1{`RANDOM}};
  _T_1718_im = _RAND_3033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3034 = {1{`RANDOM}};
  _T_1719_re = _RAND_3034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3035 = {1{`RANDOM}};
  _T_1719_im = _RAND_3035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3036 = {1{`RANDOM}};
  _T_1720_re = _RAND_3036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3037 = {1{`RANDOM}};
  _T_1720_im = _RAND_3037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3038 = {1{`RANDOM}};
  _T_1721_re = _RAND_3038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3039 = {1{`RANDOM}};
  _T_1721_im = _RAND_3039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3040 = {1{`RANDOM}};
  _T_1722_re = _RAND_3040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3041 = {1{`RANDOM}};
  _T_1722_im = _RAND_3041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3042 = {1{`RANDOM}};
  _T_1725_re = _RAND_3042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3043 = {1{`RANDOM}};
  _T_1725_im = _RAND_3043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3044 = {1{`RANDOM}};
  _T_1726_re = _RAND_3044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3045 = {1{`RANDOM}};
  _T_1726_im = _RAND_3045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3046 = {1{`RANDOM}};
  _T_1727_re = _RAND_3046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3047 = {1{`RANDOM}};
  _T_1727_im = _RAND_3047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3048 = {1{`RANDOM}};
  _T_1728_re = _RAND_3048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3049 = {1{`RANDOM}};
  _T_1728_im = _RAND_3049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3050 = {1{`RANDOM}};
  _T_1734_re = _RAND_3050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3051 = {1{`RANDOM}};
  _T_1734_im = _RAND_3051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3052 = {1{`RANDOM}};
  _T_1735_re = _RAND_3052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3053 = {1{`RANDOM}};
  _T_1735_im = _RAND_3053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3054 = {1{`RANDOM}};
  _T_1736_re = _RAND_3054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3055 = {1{`RANDOM}};
  _T_1736_im = _RAND_3055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3056 = {1{`RANDOM}};
  _T_1737_re = _RAND_3056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3057 = {1{`RANDOM}};
  _T_1737_im = _RAND_3057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3058 = {1{`RANDOM}};
  _T_1740_re = _RAND_3058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3059 = {1{`RANDOM}};
  _T_1740_im = _RAND_3059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3060 = {1{`RANDOM}};
  _T_1741_re = _RAND_3060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3061 = {1{`RANDOM}};
  _T_1741_im = _RAND_3061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3062 = {1{`RANDOM}};
  _T_1747_re = _RAND_3062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3063 = {1{`RANDOM}};
  _T_1747_im = _RAND_3063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3064 = {1{`RANDOM}};
  _T_1748_re = _RAND_3064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3065 = {1{`RANDOM}};
  _T_1748_im = _RAND_3065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3066 = {1{`RANDOM}};
  _T_1751_re = _RAND_3066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3067 = {1{`RANDOM}};
  _T_1751_im = _RAND_3067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3068 = {1{`RANDOM}};
  out1D1_re = _RAND_3068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3069 = {1{`RANDOM}};
  out1D1_im = _RAND_3069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3070 = {1{`RANDOM}};
  _T_1752_re = _RAND_3070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3071 = {1{`RANDOM}};
  _T_1752_im = _RAND_3071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3072 = {1{`RANDOM}};
  _T_1753_re = _RAND_3072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3073 = {1{`RANDOM}};
  _T_1753_im = _RAND_3073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 10'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    cntD1 <= cnt;
    _T_161_re <= io_dIn_re;
    _T_161_im <= io_dIn_im;
    _T_162_re <= _T_161_re;
    _T_162_im <= _T_161_im;
    _T_163_re <= _T_162_re;
    _T_163_im <= _T_162_im;
    _T_164_re <= _T_163_re;
    _T_164_im <= _T_163_im;
    _T_165_re <= _T_164_re;
    _T_165_im <= _T_164_im;
    _T_166_re <= _T_165_re;
    _T_166_im <= _T_165_im;
    _T_167_re <= _T_166_re;
    _T_167_im <= _T_166_im;
    _T_168_re <= _T_167_re;
    _T_168_im <= _T_167_im;
    _T_169_re <= _T_168_re;
    _T_169_im <= _T_168_im;
    _T_170_re <= _T_169_re;
    _T_170_im <= _T_169_im;
    _T_171_re <= _T_170_re;
    _T_171_im <= _T_170_im;
    _T_172_re <= _T_171_re;
    _T_172_im <= _T_171_im;
    _T_173_re <= _T_172_re;
    _T_173_im <= _T_172_im;
    _T_174_re <= _T_173_re;
    _T_174_im <= _T_173_im;
    _T_175_re <= _T_174_re;
    _T_175_im <= _T_174_im;
    _T_176_re <= _T_175_re;
    _T_176_im <= _T_175_im;
    _T_177_re <= _T_176_re;
    _T_177_im <= _T_176_im;
    _T_178_re <= _T_177_re;
    _T_178_im <= _T_177_im;
    _T_179_re <= _T_178_re;
    _T_179_im <= _T_178_im;
    _T_180_re <= _T_179_re;
    _T_180_im <= _T_179_im;
    _T_181_re <= _T_180_re;
    _T_181_im <= _T_180_im;
    _T_182_re <= _T_181_re;
    _T_182_im <= _T_181_im;
    _T_183_re <= _T_182_re;
    _T_183_im <= _T_182_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_325_re <= _T_324_re;
    _T_325_im <= _T_324_im;
    _T_326_re <= _T_325_re;
    _T_326_im <= _T_325_im;
    _T_327_re <= _T_326_re;
    _T_327_im <= _T_326_im;
    _T_328_re <= _T_327_re;
    _T_328_im <= _T_327_im;
    _T_329_re <= _T_328_re;
    _T_329_im <= _T_328_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_393_re <= _T_392_re;
    _T_393_im <= _T_392_im;
    _T_394_re <= _T_393_re;
    _T_394_im <= _T_393_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_402_re <= _T_401_re;
    _T_402_im <= _T_401_im;
    _T_403_re <= _T_402_re;
    _T_403_im <= _T_402_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_406_re <= _T_405_re;
    _T_406_im <= _T_405_im;
    _T_407_re <= _T_406_re;
    _T_407_im <= _T_406_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_409_re <= _T_408_re;
    _T_409_im <= _T_408_im;
    _T_410_re <= _T_409_re;
    _T_410_im <= _T_409_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_533_re <= _T_532_re;
    _T_533_im <= _T_532_im;
    _T_534_re <= _T_533_re;
    _T_534_im <= _T_533_im;
    _T_535_re <= _T_534_re;
    _T_535_im <= _T_534_im;
    _T_536_re <= _T_535_re;
    _T_536_im <= _T_535_im;
    _T_537_re <= _T_536_re;
    _T_537_im <= _T_536_im;
    _T_538_re <= _T_537_re;
    _T_538_im <= _T_537_im;
    _T_539_re <= _T_538_re;
    _T_539_im <= _T_538_im;
    _T_540_re <= _T_539_re;
    _T_540_im <= _T_539_im;
    _T_541_re <= _T_540_re;
    _T_541_im <= _T_540_im;
    _T_542_re <= _T_541_re;
    _T_542_im <= _T_541_im;
    _T_543_re <= _T_542_re;
    _T_543_im <= _T_542_im;
    _T_544_re <= _T_543_re;
    _T_544_im <= _T_543_im;
    _T_545_re <= _T_544_re;
    _T_545_im <= _T_544_im;
    _T_546_re <= _T_545_re;
    _T_546_im <= _T_545_im;
    _T_547_re <= _T_546_re;
    _T_547_im <= _T_546_im;
    _T_548_re <= _T_547_re;
    _T_548_im <= _T_547_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_663_re <= _T_662_re;
    _T_663_im <= _T_662_im;
    _T_664_re <= _T_663_re;
    _T_664_im <= _T_663_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_671_re <= _T_670_re;
    _T_671_im <= _T_670_im;
    _T_672_re <= _T_671_re;
    _T_672_im <= _T_671_im;
    _T_675_re <= Butterfly_io_out2_re;
    _T_675_im <= Butterfly_io_out2_im;
    _T_676_re <= _T_675_re;
    _T_676_im <= _T_675_im;
    _T_677_re <= _T_676_re;
    _T_677_im <= _T_676_im;
    _T_678_re <= _T_677_re;
    _T_678_im <= _T_677_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_728_re <= _T_727_re;
    _T_728_im <= _T_727_im;
    _T_729_re <= _T_728_re;
    _T_729_im <= _T_728_im;
    _T_730_re <= _T_729_re;
    _T_730_im <= _T_729_im;
    _T_731_re <= _T_730_re;
    _T_731_im <= _T_730_im;
    _T_732_re <= _T_731_re;
    _T_732_im <= _T_731_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_736_re <= _T_735_re;
    _T_736_im <= _T_735_im;
    _T_737_re <= _T_736_re;
    _T_737_im <= _T_736_im;
    _T_738_re <= _T_737_re;
    _T_738_im <= _T_737_im;
    _T_739_re <= _T_738_re;
    _T_739_im <= _T_738_im;
    _T_740_re <= _T_739_re;
    _T_740_im <= _T_739_im;
    _T_741_re <= _T_740_re;
    _T_741_im <= _T_740_im;
    _T_742_re <= _T_741_re;
    _T_742_im <= _T_741_im;
    _T_743_re <= _T_742_re;
    _T_743_im <= _T_742_im;
    _T_744_re <= _T_743_re;
    _T_744_im <= _T_743_im;
    _T_745_re <= _T_744_re;
    _T_745_im <= _T_744_im;
    _T_746_re <= _T_745_re;
    _T_746_im <= _T_745_im;
    _T_747_re <= _T_746_re;
    _T_747_im <= _T_746_im;
    _T_748_re <= _T_747_re;
    _T_748_im <= _T_747_im;
    _T_749_re <= _T_748_re;
    _T_749_im <= _T_748_im;
    _T_750_re <= _T_749_re;
    _T_750_im <= _T_749_im;
    _T_751_re <= _T_750_re;
    _T_751_im <= _T_750_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_796_re <= _T_795_re;
    _T_796_im <= _T_795_im;
    _T_797_re <= _T_796_re;
    _T_797_im <= _T_796_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_808_re <= _T_807_re;
    _T_808_im <= _T_807_im;
    _T_809_re <= _T_808_re;
    _T_809_im <= _T_808_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_811_re <= _T_810_re;
    _T_811_im <= _T_810_im;
    _T_812_re <= _T_811_re;
    _T_812_im <= _T_811_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_815_re <= _T_814_re;
    _T_815_im <= _T_814_im;
    _T_816_re <= _T_815_re;
    _T_816_im <= _T_815_im;
    _T_817_re <= _T_816_re;
    _T_817_im <= _T_816_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_829_re <= _T_828_re;
    _T_829_im <= _T_828_im;
    _T_830_re <= _T_829_re;
    _T_830_im <= _T_829_im;
    _T_831_re <= _T_830_re;
    _T_831_im <= _T_830_im;
    _T_832_re <= _T_831_re;
    _T_832_im <= _T_831_im;
    _T_833_re <= _T_832_re;
    _T_833_im <= _T_832_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_841_re <= _T_840_re;
    _T_841_im <= _T_840_im;
    _T_842_re <= _T_841_re;
    _T_842_im <= _T_841_im;
    _T_843_re <= _T_842_re;
    _T_843_im <= _T_842_im;
    _T_844_re <= _T_843_re;
    _T_844_im <= _T_843_im;
    _T_845_re <= _T_844_re;
    _T_845_im <= _T_844_im;
    _T_846_re <= _T_845_re;
    _T_846_im <= _T_845_im;
    _T_847_re <= _T_846_re;
    _T_847_im <= _T_846_im;
    _T_848_re <= _T_847_re;
    _T_848_im <= _T_847_im;
    _T_849_re <= _T_848_re;
    _T_849_im <= _T_848_im;
    _T_850_re <= _T_849_re;
    _T_850_im <= _T_849_im;
    _T_851_re <= _T_850_re;
    _T_851_im <= _T_850_im;
    _T_852_re <= _T_851_re;
    _T_852_im <= _T_851_im;
    _T_853_re <= _T_852_re;
    _T_853_im <= _T_852_im;
    _T_854_re <= _T_853_re;
    _T_854_im <= _T_853_im;
    _T_855_re <= _T_854_re;
    _T_855_im <= _T_854_im;
    _T_856_re <= _T_855_re;
    _T_856_im <= _T_855_im;
    _T_857_re <= _T_856_re;
    _T_857_im <= _T_856_im;
    _T_858_re <= _T_857_re;
    _T_858_im <= _T_857_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_865_re <= _T_864_re;
    _T_865_im <= _T_864_im;
    _T_866_re <= _T_865_re;
    _T_866_im <= _T_865_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_881_re <= _T_880_re;
    _T_881_im <= _T_880_im;
    _T_882_re <= _T_881_re;
    _T_882_im <= _T_881_im;
    _T_883_re <= _T_882_re;
    _T_883_im <= _T_882_im;
    _T_884_re <= _T_883_re;
    _T_884_im <= _T_883_im;
    _T_885_re <= _T_884_re;
    _T_885_im <= _T_884_im;
    _T_886_re <= _T_885_re;
    _T_886_im <= _T_885_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_890_re <= _T_889_re;
    _T_890_im <= _T_889_im;
    _T_891_re <= _T_890_re;
    _T_891_im <= _T_890_im;
    _T_892_re <= _T_891_re;
    _T_892_im <= _T_891_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_898_re <= _T_897_re;
    _T_898_im <= _T_897_im;
    _T_899_re <= _T_898_re;
    _T_899_im <= _T_898_im;
    _T_900_re <= _T_899_re;
    _T_900_im <= _T_899_im;
    _T_901_re <= _T_900_re;
    _T_901_im <= _T_900_im;
    _T_902_re <= _T_901_re;
    _T_902_im <= _T_901_im;
    _T_903_re <= _T_902_re;
    _T_903_im <= _T_902_im;
    _T_904_re <= _T_903_re;
    _T_904_im <= _T_903_im;
    _T_905_re <= _T_904_re;
    _T_905_im <= _T_904_im;
    _T_906_re <= _T_905_re;
    _T_906_im <= _T_905_im;
    _T_907_re <= _T_906_re;
    _T_907_im <= _T_906_im;
    _T_908_re <= _T_907_re;
    _T_908_im <= _T_907_im;
    _T_909_re <= _T_908_re;
    _T_909_im <= _T_908_im;
    _T_910_re <= _T_909_re;
    _T_910_im <= _T_909_im;
    _T_911_re <= _T_910_re;
    _T_911_im <= _T_910_im;
    _T_912_re <= _T_911_re;
    _T_912_im <= _T_911_im;
    _T_913_re <= _T_912_re;
    _T_913_im <= _T_912_im;
    _T_914_re <= _T_913_re;
    _T_914_im <= _T_913_im;
    _T_915_re <= _T_914_re;
    _T_915_im <= _T_914_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_922_re <= _T_921_re;
    _T_922_im <= _T_921_im;
    _T_923_re <= _T_922_re;
    _T_923_im <= _T_922_im;
    _T_924_re <= _T_923_re;
    _T_924_im <= _T_923_im;
    _T_925_re <= _T_924_re;
    _T_925_im <= _T_924_im;
    _T_926_re <= _T_925_re;
    _T_926_im <= _T_925_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_928_re <= _T_927_re;
    _T_928_im <= _T_927_im;
    _T_929_re <= _T_928_re;
    _T_929_im <= _T_928_im;
    _T_930_re <= _T_929_re;
    _T_930_im <= _T_929_im;
    _T_936_re <= Switch_io_out1_re;
    _T_936_im <= Switch_io_out1_im;
    _T_937_re <= _T_936_re;
    _T_937_im <= _T_936_im;
    _T_938_re <= _T_937_re;
    _T_938_im <= _T_937_im;
    _T_939_re <= _T_938_re;
    _T_939_im <= _T_938_im;
    _T_940_re <= _T_939_re;
    _T_940_im <= _T_939_im;
    _T_941_re <= _T_940_re;
    _T_941_im <= _T_940_im;
    _T_942_re <= _T_941_re;
    _T_942_im <= _T_941_im;
    _T_943_re <= _T_942_re;
    _T_943_im <= _T_942_im;
    _T_944_re <= _T_943_re;
    _T_944_im <= _T_943_im;
    _T_945_re <= _T_944_re;
    _T_945_im <= _T_944_im;
    _T_946_re <= _T_945_re;
    _T_946_im <= _T_945_im;
    _T_947_re <= _T_946_re;
    _T_947_im <= _T_946_im;
    _T_948_re <= _T_947_re;
    _T_948_im <= _T_947_im;
    _T_949_re <= _T_948_re;
    _T_949_im <= _T_948_im;
    _T_950_re <= _T_949_re;
    _T_950_im <= _T_949_im;
    _T_951_re <= _T_950_re;
    _T_951_im <= _T_950_im;
    _T_952_re <= _T_951_re;
    _T_952_im <= _T_951_im;
    _T_953_re <= _T_952_re;
    _T_953_im <= _T_952_im;
    _T_954_re <= _T_953_re;
    _T_954_im <= _T_953_im;
    _T_955_re <= _T_954_re;
    _T_955_im <= _T_954_im;
    _T_956_re <= _T_955_re;
    _T_956_im <= _T_955_im;
    _T_957_re <= _T_956_re;
    _T_957_im <= _T_956_im;
    _T_958_re <= _T_957_re;
    _T_958_im <= _T_957_im;
    _T_959_re <= _T_958_re;
    _T_959_im <= _T_958_im;
    _T_960_re <= _T_959_re;
    _T_960_im <= _T_959_im;
    _T_961_re <= _T_960_re;
    _T_961_im <= _T_960_im;
    _T_962_re <= _T_961_re;
    _T_962_im <= _T_961_im;
    _T_963_re <= _T_962_re;
    _T_963_im <= _T_962_im;
    _T_964_re <= _T_963_re;
    _T_964_im <= _T_963_im;
    _T_965_re <= _T_964_re;
    _T_965_im <= _T_964_im;
    _T_966_re <= _T_965_re;
    _T_966_im <= _T_965_im;
    _T_967_re <= _T_966_re;
    _T_967_im <= _T_966_im;
    _T_968_re <= _T_967_re;
    _T_968_im <= _T_967_im;
    _T_969_re <= _T_968_re;
    _T_969_im <= _T_968_im;
    _T_970_re <= _T_969_re;
    _T_970_im <= _T_969_im;
    _T_971_re <= _T_970_re;
    _T_971_im <= _T_970_im;
    _T_972_re <= _T_971_re;
    _T_972_im <= _T_971_im;
    _T_973_re <= _T_972_re;
    _T_973_im <= _T_972_im;
    _T_974_re <= _T_973_re;
    _T_974_im <= _T_973_im;
    _T_975_re <= _T_974_re;
    _T_975_im <= _T_974_im;
    _T_976_re <= _T_975_re;
    _T_976_im <= _T_975_im;
    _T_977_re <= _T_976_re;
    _T_977_im <= _T_976_im;
    _T_978_re <= _T_977_re;
    _T_978_im <= _T_977_im;
    _T_979_re <= _T_978_re;
    _T_979_im <= _T_978_im;
    _T_980_re <= _T_979_re;
    _T_980_im <= _T_979_im;
    _T_981_re <= _T_980_re;
    _T_981_im <= _T_980_im;
    _T_982_re <= _T_981_re;
    _T_982_im <= _T_981_im;
    _T_983_re <= _T_982_re;
    _T_983_im <= _T_982_im;
    _T_984_re <= _T_983_re;
    _T_984_im <= _T_983_im;
    _T_985_re <= _T_984_re;
    _T_985_im <= _T_984_im;
    _T_986_re <= _T_985_re;
    _T_986_im <= _T_985_im;
    _T_987_re <= _T_986_re;
    _T_987_im <= _T_986_im;
    _T_988_re <= _T_987_re;
    _T_988_im <= _T_987_im;
    _T_989_re <= _T_988_re;
    _T_989_im <= _T_988_im;
    _T_990_re <= _T_989_re;
    _T_990_im <= _T_989_im;
    _T_991_re <= _T_990_re;
    _T_991_im <= _T_990_im;
    _T_992_re <= _T_991_re;
    _T_992_im <= _T_991_im;
    _T_993_re <= _T_992_re;
    _T_993_im <= _T_992_im;
    _T_994_re <= _T_993_re;
    _T_994_im <= _T_993_im;
    _T_995_re <= _T_994_re;
    _T_995_im <= _T_994_im;
    _T_996_re <= _T_995_re;
    _T_996_im <= _T_995_im;
    _T_997_re <= _T_996_re;
    _T_997_im <= _T_996_im;
    _T_998_re <= _T_997_re;
    _T_998_im <= _T_997_im;
    _T_999_re <= _T_998_re;
    _T_999_im <= _T_998_im;
    _T_1000_re <= _T_999_re;
    _T_1000_im <= _T_999_im;
    _T_1001_re <= _T_1000_re;
    _T_1001_im <= _T_1000_im;
    _T_1002_re <= _T_1001_re;
    _T_1002_im <= _T_1001_im;
    _T_1003_re <= _T_1002_re;
    _T_1003_im <= _T_1002_im;
    _T_1004_re <= _T_1003_re;
    _T_1004_im <= _T_1003_im;
    _T_1005_re <= _T_1004_re;
    _T_1005_im <= _T_1004_im;
    _T_1006_re <= _T_1005_re;
    _T_1006_im <= _T_1005_im;
    _T_1007_re <= _T_1006_re;
    _T_1007_im <= _T_1006_im;
    _T_1008_re <= _T_1007_re;
    _T_1008_im <= _T_1007_im;
    _T_1009_re <= _T_1008_re;
    _T_1009_im <= _T_1008_im;
    _T_1010_re <= _T_1009_re;
    _T_1010_im <= _T_1009_im;
    _T_1011_re <= _T_1010_re;
    _T_1011_im <= _T_1010_im;
    _T_1012_re <= _T_1011_re;
    _T_1012_im <= _T_1011_im;
    _T_1013_re <= _T_1012_re;
    _T_1013_im <= _T_1012_im;
    _T_1014_re <= _T_1013_re;
    _T_1014_im <= _T_1013_im;
    _T_1015_re <= _T_1014_re;
    _T_1015_im <= _T_1014_im;
    _T_1016_re <= _T_1015_re;
    _T_1016_im <= _T_1015_im;
    _T_1017_re <= _T_1016_re;
    _T_1017_im <= _T_1016_im;
    _T_1018_re <= _T_1017_re;
    _T_1018_im <= _T_1017_im;
    _T_1019_re <= _T_1018_re;
    _T_1019_im <= _T_1018_im;
    _T_1020_re <= _T_1019_re;
    _T_1020_im <= _T_1019_im;
    _T_1021_re <= _T_1020_re;
    _T_1021_im <= _T_1020_im;
    _T_1022_re <= _T_1021_re;
    _T_1022_im <= _T_1021_im;
    _T_1023_re <= _T_1022_re;
    _T_1023_im <= _T_1022_im;
    _T_1024_re <= _T_1023_re;
    _T_1024_im <= _T_1023_im;
    _T_1025_re <= _T_1024_re;
    _T_1025_im <= _T_1024_im;
    _T_1026_re <= _T_1025_re;
    _T_1026_im <= _T_1025_im;
    _T_1027_re <= _T_1026_re;
    _T_1027_im <= _T_1026_im;
    _T_1028_re <= _T_1027_re;
    _T_1028_im <= _T_1027_im;
    _T_1029_re <= _T_1028_re;
    _T_1029_im <= _T_1028_im;
    _T_1030_re <= _T_1029_re;
    _T_1030_im <= _T_1029_im;
    _T_1031_re <= _T_1030_re;
    _T_1031_im <= _T_1030_im;
    _T_1032_re <= _T_1031_re;
    _T_1032_im <= _T_1031_im;
    _T_1033_re <= _T_1032_re;
    _T_1033_im <= _T_1032_im;
    _T_1034_re <= _T_1033_re;
    _T_1034_im <= _T_1033_im;
    _T_1035_re <= _T_1034_re;
    _T_1035_im <= _T_1034_im;
    _T_1036_re <= _T_1035_re;
    _T_1036_im <= _T_1035_im;
    _T_1037_re <= _T_1036_re;
    _T_1037_im <= _T_1036_im;
    _T_1038_re <= _T_1037_re;
    _T_1038_im <= _T_1037_im;
    _T_1039_re <= _T_1038_re;
    _T_1039_im <= _T_1038_im;
    _T_1040_re <= _T_1039_re;
    _T_1040_im <= _T_1039_im;
    _T_1041_re <= _T_1040_re;
    _T_1041_im <= _T_1040_im;
    _T_1042_re <= _T_1041_re;
    _T_1042_im <= _T_1041_im;
    _T_1043_re <= _T_1042_re;
    _T_1043_im <= _T_1042_im;
    _T_1044_re <= _T_1043_re;
    _T_1044_im <= _T_1043_im;
    _T_1045_re <= _T_1044_re;
    _T_1045_im <= _T_1044_im;
    _T_1046_re <= _T_1045_re;
    _T_1046_im <= _T_1045_im;
    _T_1047_re <= _T_1046_re;
    _T_1047_im <= _T_1046_im;
    _T_1048_re <= _T_1047_re;
    _T_1048_im <= _T_1047_im;
    _T_1049_re <= _T_1048_re;
    _T_1049_im <= _T_1048_im;
    _T_1050_re <= _T_1049_re;
    _T_1050_im <= _T_1049_im;
    _T_1051_re <= _T_1050_re;
    _T_1051_im <= _T_1050_im;
    _T_1052_re <= _T_1051_re;
    _T_1052_im <= _T_1051_im;
    _T_1053_re <= _T_1052_re;
    _T_1053_im <= _T_1052_im;
    _T_1054_re <= _T_1053_re;
    _T_1054_im <= _T_1053_im;
    _T_1055_re <= _T_1054_re;
    _T_1055_im <= _T_1054_im;
    _T_1056_re <= _T_1055_re;
    _T_1056_im <= _T_1055_im;
    _T_1057_re <= _T_1056_re;
    _T_1057_im <= _T_1056_im;
    _T_1058_re <= _T_1057_re;
    _T_1058_im <= _T_1057_im;
    _T_1059_re <= _T_1058_re;
    _T_1059_im <= _T_1058_im;
    _T_1060_re <= _T_1059_re;
    _T_1060_im <= _T_1059_im;
    _T_1061_re <= _T_1060_re;
    _T_1061_im <= _T_1060_im;
    _T_1062_re <= _T_1061_re;
    _T_1062_im <= _T_1061_im;
    _T_1063_re <= _T_1062_re;
    _T_1063_im <= _T_1062_im;
    _T_1064_re <= _T_1063_re;
    _T_1064_im <= _T_1063_im;
    _T_1065_re <= _T_1064_re;
    _T_1065_im <= _T_1064_im;
    _T_1066_re <= _T_1065_re;
    _T_1066_im <= _T_1065_im;
    _T_1067_re <= _T_1066_re;
    _T_1067_im <= _T_1066_im;
    _T_1068_re <= _T_1067_re;
    _T_1068_im <= _T_1067_im;
    _T_1069_re <= _T_1068_re;
    _T_1069_im <= _T_1068_im;
    _T_1070_re <= _T_1069_re;
    _T_1070_im <= _T_1069_im;
    _T_1071_re <= _T_1070_re;
    _T_1071_im <= _T_1070_im;
    _T_1072_re <= _T_1071_re;
    _T_1072_im <= _T_1071_im;
    _T_1073_re <= _T_1072_re;
    _T_1073_im <= _T_1072_im;
    _T_1074_re <= _T_1073_re;
    _T_1074_im <= _T_1073_im;
    _T_1075_re <= _T_1074_re;
    _T_1075_im <= _T_1074_im;
    _T_1076_re <= _T_1075_re;
    _T_1076_im <= _T_1075_im;
    _T_1077_re <= _T_1076_re;
    _T_1077_im <= _T_1076_im;
    _T_1078_re <= _T_1077_re;
    _T_1078_im <= _T_1077_im;
    _T_1079_re <= _T_1078_re;
    _T_1079_im <= _T_1078_im;
    _T_1080_re <= _T_1079_re;
    _T_1080_im <= _T_1079_im;
    _T_1081_re <= _T_1080_re;
    _T_1081_im <= _T_1080_im;
    _T_1082_re <= _T_1081_re;
    _T_1082_im <= _T_1081_im;
    _T_1083_re <= _T_1082_re;
    _T_1083_im <= _T_1082_im;
    _T_1084_re <= _T_1083_re;
    _T_1084_im <= _T_1083_im;
    _T_1085_re <= _T_1084_re;
    _T_1085_im <= _T_1084_im;
    _T_1086_re <= _T_1085_re;
    _T_1086_im <= _T_1085_im;
    _T_1087_re <= _T_1086_re;
    _T_1087_im <= _T_1086_im;
    _T_1088_re <= _T_1087_re;
    _T_1088_im <= _T_1087_im;
    _T_1089_re <= _T_1088_re;
    _T_1089_im <= _T_1088_im;
    _T_1090_re <= _T_1089_re;
    _T_1090_im <= _T_1089_im;
    _T_1091_re <= _T_1090_re;
    _T_1091_im <= _T_1090_im;
    _T_1092_re <= _T_1091_re;
    _T_1092_im <= _T_1091_im;
    _T_1093_re <= _T_1092_re;
    _T_1093_im <= _T_1092_im;
    _T_1094_re <= _T_1093_re;
    _T_1094_im <= _T_1093_im;
    _T_1095_re <= _T_1094_re;
    _T_1095_im <= _T_1094_im;
    _T_1096_re <= _T_1095_re;
    _T_1096_im <= _T_1095_im;
    _T_1097_re <= _T_1096_re;
    _T_1097_im <= _T_1096_im;
    _T_1098_re <= _T_1097_re;
    _T_1098_im <= _T_1097_im;
    _T_1099_re <= _T_1098_re;
    _T_1099_im <= _T_1098_im;
    _T_1100_re <= _T_1099_re;
    _T_1100_im <= _T_1099_im;
    _T_1101_re <= _T_1100_re;
    _T_1101_im <= _T_1100_im;
    _T_1102_re <= _T_1101_re;
    _T_1102_im <= _T_1101_im;
    _T_1103_re <= _T_1102_re;
    _T_1103_im <= _T_1102_im;
    _T_1104_re <= _T_1103_re;
    _T_1104_im <= _T_1103_im;
    _T_1105_re <= _T_1104_re;
    _T_1105_im <= _T_1104_im;
    _T_1106_re <= _T_1105_re;
    _T_1106_im <= _T_1105_im;
    _T_1107_re <= _T_1106_re;
    _T_1107_im <= _T_1106_im;
    _T_1108_re <= _T_1107_re;
    _T_1108_im <= _T_1107_im;
    _T_1109_re <= _T_1108_re;
    _T_1109_im <= _T_1108_im;
    _T_1110_re <= _T_1109_re;
    _T_1110_im <= _T_1109_im;
    _T_1111_re <= _T_1110_re;
    _T_1111_im <= _T_1110_im;
    _T_1112_re <= _T_1111_re;
    _T_1112_im <= _T_1111_im;
    _T_1113_re <= _T_1112_re;
    _T_1113_im <= _T_1112_im;
    _T_1114_re <= _T_1113_re;
    _T_1114_im <= _T_1113_im;
    _T_1115_re <= _T_1114_re;
    _T_1115_im <= _T_1114_im;
    _T_1116_re <= _T_1115_re;
    _T_1116_im <= _T_1115_im;
    _T_1117_re <= _T_1116_re;
    _T_1117_im <= _T_1116_im;
    _T_1118_re <= _T_1117_re;
    _T_1118_im <= _T_1117_im;
    _T_1119_re <= _T_1118_re;
    _T_1119_im <= _T_1118_im;
    _T_1120_re <= _T_1119_re;
    _T_1120_im <= _T_1119_im;
    _T_1121_re <= _T_1120_re;
    _T_1121_im <= _T_1120_im;
    _T_1122_re <= _T_1121_re;
    _T_1122_im <= _T_1121_im;
    _T_1123_re <= _T_1122_re;
    _T_1123_im <= _T_1122_im;
    _T_1124_re <= _T_1123_re;
    _T_1124_im <= _T_1123_im;
    _T_1125_re <= _T_1124_re;
    _T_1125_im <= _T_1124_im;
    _T_1126_re <= _T_1125_re;
    _T_1126_im <= _T_1125_im;
    _T_1127_re <= _T_1126_re;
    _T_1127_im <= _T_1126_im;
    _T_1128_re <= _T_1127_re;
    _T_1128_im <= _T_1127_im;
    _T_1129_re <= _T_1128_re;
    _T_1129_im <= _T_1128_im;
    _T_1130_re <= _T_1129_re;
    _T_1130_im <= _T_1129_im;
    _T_1131_re <= _T_1130_re;
    _T_1131_im <= _T_1130_im;
    _T_1132_re <= _T_1131_re;
    _T_1132_im <= _T_1131_im;
    _T_1133_re <= _T_1132_re;
    _T_1133_im <= _T_1132_im;
    _T_1134_re <= _T_1133_re;
    _T_1134_im <= _T_1133_im;
    _T_1135_re <= _T_1134_re;
    _T_1135_im <= _T_1134_im;
    _T_1136_re <= _T_1135_re;
    _T_1136_im <= _T_1135_im;
    _T_1137_re <= _T_1136_re;
    _T_1137_im <= _T_1136_im;
    _T_1138_re <= _T_1137_re;
    _T_1138_im <= _T_1137_im;
    _T_1139_re <= _T_1138_re;
    _T_1139_im <= _T_1138_im;
    _T_1140_re <= _T_1139_re;
    _T_1140_im <= _T_1139_im;
    _T_1141_re <= _T_1140_re;
    _T_1141_im <= _T_1140_im;
    _T_1142_re <= _T_1141_re;
    _T_1142_im <= _T_1141_im;
    _T_1143_re <= _T_1142_re;
    _T_1143_im <= _T_1142_im;
    _T_1144_re <= _T_1143_re;
    _T_1144_im <= _T_1143_im;
    _T_1145_re <= _T_1144_re;
    _T_1145_im <= _T_1144_im;
    _T_1146_re <= _T_1145_re;
    _T_1146_im <= _T_1145_im;
    _T_1147_re <= _T_1146_re;
    _T_1147_im <= _T_1146_im;
    _T_1148_re <= _T_1147_re;
    _T_1148_im <= _T_1147_im;
    _T_1149_re <= _T_1148_re;
    _T_1149_im <= _T_1148_im;
    _T_1150_re <= _T_1149_re;
    _T_1150_im <= _T_1149_im;
    _T_1151_re <= _T_1150_re;
    _T_1151_im <= _T_1150_im;
    _T_1152_re <= _T_1151_re;
    _T_1152_im <= _T_1151_im;
    _T_1153_re <= _T_1152_re;
    _T_1153_im <= _T_1152_im;
    _T_1154_re <= _T_1153_re;
    _T_1154_im <= _T_1153_im;
    _T_1155_re <= _T_1154_re;
    _T_1155_im <= _T_1154_im;
    _T_1156_re <= _T_1155_re;
    _T_1156_im <= _T_1155_im;
    _T_1157_re <= _T_1156_re;
    _T_1157_im <= _T_1156_im;
    _T_1158_re <= _T_1157_re;
    _T_1158_im <= _T_1157_im;
    _T_1159_re <= _T_1158_re;
    _T_1159_im <= _T_1158_im;
    _T_1160_re <= _T_1159_re;
    _T_1160_im <= _T_1159_im;
    _T_1161_re <= _T_1160_re;
    _T_1161_im <= _T_1160_im;
    _T_1162_re <= _T_1161_re;
    _T_1162_im <= _T_1161_im;
    _T_1163_re <= _T_1162_re;
    _T_1163_im <= _T_1162_im;
    _T_1164_re <= _T_1163_re;
    _T_1164_im <= _T_1163_im;
    _T_1165_re <= _T_1164_re;
    _T_1165_im <= _T_1164_im;
    _T_1166_re <= _T_1165_re;
    _T_1166_im <= _T_1165_im;
    _T_1167_re <= _T_1166_re;
    _T_1167_im <= _T_1166_im;
    _T_1168_re <= _T_1167_re;
    _T_1168_im <= _T_1167_im;
    _T_1169_re <= _T_1168_re;
    _T_1169_im <= _T_1168_im;
    _T_1170_re <= _T_1169_re;
    _T_1170_im <= _T_1169_im;
    _T_1171_re <= _T_1170_re;
    _T_1171_im <= _T_1170_im;
    _T_1172_re <= _T_1171_re;
    _T_1172_im <= _T_1171_im;
    _T_1173_re <= _T_1172_re;
    _T_1173_im <= _T_1172_im;
    _T_1174_re <= _T_1173_re;
    _T_1174_im <= _T_1173_im;
    _T_1175_re <= _T_1174_re;
    _T_1175_im <= _T_1174_im;
    _T_1176_re <= _T_1175_re;
    _T_1176_im <= _T_1175_im;
    _T_1177_re <= _T_1176_re;
    _T_1177_im <= _T_1176_im;
    _T_1178_re <= _T_1177_re;
    _T_1178_im <= _T_1177_im;
    _T_1179_re <= _T_1178_re;
    _T_1179_im <= _T_1178_im;
    _T_1180_re <= _T_1179_re;
    _T_1180_im <= _T_1179_im;
    _T_1181_re <= _T_1180_re;
    _T_1181_im <= _T_1180_im;
    _T_1182_re <= _T_1181_re;
    _T_1182_im <= _T_1181_im;
    _T_1183_re <= _T_1182_re;
    _T_1183_im <= _T_1182_im;
    _T_1184_re <= _T_1183_re;
    _T_1184_im <= _T_1183_im;
    _T_1185_re <= _T_1184_re;
    _T_1185_im <= _T_1184_im;
    _T_1186_re <= _T_1185_re;
    _T_1186_im <= _T_1185_im;
    _T_1187_re <= _T_1186_re;
    _T_1187_im <= _T_1186_im;
    _T_1188_re <= _T_1187_re;
    _T_1188_im <= _T_1187_im;
    _T_1189_re <= _T_1188_re;
    _T_1189_im <= _T_1188_im;
    _T_1190_re <= _T_1189_re;
    _T_1190_im <= _T_1189_im;
    _T_1191_re <= _T_1190_re;
    _T_1191_im <= _T_1190_im;
    _T_1194_re <= Butterfly_1_io_out2_re;
    _T_1194_im <= Butterfly_1_io_out2_im;
    _T_1195_re <= _T_1194_re;
    _T_1195_im <= _T_1194_im;
    _T_1196_re <= _T_1195_re;
    _T_1196_im <= _T_1195_im;
    _T_1197_re <= _T_1196_re;
    _T_1197_im <= _T_1196_im;
    _T_1198_re <= _T_1197_re;
    _T_1198_im <= _T_1197_im;
    _T_1199_re <= _T_1198_re;
    _T_1199_im <= _T_1198_im;
    _T_1200_re <= _T_1199_re;
    _T_1200_im <= _T_1199_im;
    _T_1201_re <= _T_1200_re;
    _T_1201_im <= _T_1200_im;
    _T_1202_re <= _T_1201_re;
    _T_1202_im <= _T_1201_im;
    _T_1203_re <= _T_1202_re;
    _T_1203_im <= _T_1202_im;
    _T_1204_re <= _T_1203_re;
    _T_1204_im <= _T_1203_im;
    _T_1205_re <= _T_1204_re;
    _T_1205_im <= _T_1204_im;
    _T_1206_re <= _T_1205_re;
    _T_1206_im <= _T_1205_im;
    _T_1207_re <= _T_1206_re;
    _T_1207_im <= _T_1206_im;
    _T_1208_re <= _T_1207_re;
    _T_1208_im <= _T_1207_im;
    _T_1209_re <= _T_1208_re;
    _T_1209_im <= _T_1208_im;
    _T_1210_re <= _T_1209_re;
    _T_1210_im <= _T_1209_im;
    _T_1211_re <= _T_1210_re;
    _T_1211_im <= _T_1210_im;
    _T_1212_re <= _T_1211_re;
    _T_1212_im <= _T_1211_im;
    _T_1213_re <= _T_1212_re;
    _T_1213_im <= _T_1212_im;
    _T_1214_re <= _T_1213_re;
    _T_1214_im <= _T_1213_im;
    _T_1215_re <= _T_1214_re;
    _T_1215_im <= _T_1214_im;
    _T_1216_re <= _T_1215_re;
    _T_1216_im <= _T_1215_im;
    _T_1217_re <= _T_1216_re;
    _T_1217_im <= _T_1216_im;
    _T_1218_re <= _T_1217_re;
    _T_1218_im <= _T_1217_im;
    _T_1219_re <= _T_1218_re;
    _T_1219_im <= _T_1218_im;
    _T_1220_re <= _T_1219_re;
    _T_1220_im <= _T_1219_im;
    _T_1221_re <= _T_1220_re;
    _T_1221_im <= _T_1220_im;
    _T_1222_re <= _T_1221_re;
    _T_1222_im <= _T_1221_im;
    _T_1223_re <= _T_1222_re;
    _T_1223_im <= _T_1222_im;
    _T_1224_re <= _T_1223_re;
    _T_1224_im <= _T_1223_im;
    _T_1225_re <= _T_1224_re;
    _T_1225_im <= _T_1224_im;
    _T_1226_re <= _T_1225_re;
    _T_1226_im <= _T_1225_im;
    _T_1227_re <= _T_1226_re;
    _T_1227_im <= _T_1226_im;
    _T_1228_re <= _T_1227_re;
    _T_1228_im <= _T_1227_im;
    _T_1229_re <= _T_1228_re;
    _T_1229_im <= _T_1228_im;
    _T_1230_re <= _T_1229_re;
    _T_1230_im <= _T_1229_im;
    _T_1231_re <= _T_1230_re;
    _T_1231_im <= _T_1230_im;
    _T_1232_re <= _T_1231_re;
    _T_1232_im <= _T_1231_im;
    _T_1233_re <= _T_1232_re;
    _T_1233_im <= _T_1232_im;
    _T_1234_re <= _T_1233_re;
    _T_1234_im <= _T_1233_im;
    _T_1235_re <= _T_1234_re;
    _T_1235_im <= _T_1234_im;
    _T_1236_re <= _T_1235_re;
    _T_1236_im <= _T_1235_im;
    _T_1237_re <= _T_1236_re;
    _T_1237_im <= _T_1236_im;
    _T_1238_re <= _T_1237_re;
    _T_1238_im <= _T_1237_im;
    _T_1239_re <= _T_1238_re;
    _T_1239_im <= _T_1238_im;
    _T_1240_re <= _T_1239_re;
    _T_1240_im <= _T_1239_im;
    _T_1241_re <= _T_1240_re;
    _T_1241_im <= _T_1240_im;
    _T_1242_re <= _T_1241_re;
    _T_1242_im <= _T_1241_im;
    _T_1243_re <= _T_1242_re;
    _T_1243_im <= _T_1242_im;
    _T_1244_re <= _T_1243_re;
    _T_1244_im <= _T_1243_im;
    _T_1245_re <= _T_1244_re;
    _T_1245_im <= _T_1244_im;
    _T_1246_re <= _T_1245_re;
    _T_1246_im <= _T_1245_im;
    _T_1247_re <= _T_1246_re;
    _T_1247_im <= _T_1246_im;
    _T_1248_re <= _T_1247_re;
    _T_1248_im <= _T_1247_im;
    _T_1249_re <= _T_1248_re;
    _T_1249_im <= _T_1248_im;
    _T_1250_re <= _T_1249_re;
    _T_1250_im <= _T_1249_im;
    _T_1251_re <= _T_1250_re;
    _T_1251_im <= _T_1250_im;
    _T_1252_re <= _T_1251_re;
    _T_1252_im <= _T_1251_im;
    _T_1253_re <= _T_1252_re;
    _T_1253_im <= _T_1252_im;
    _T_1254_re <= _T_1253_re;
    _T_1254_im <= _T_1253_im;
    _T_1255_re <= _T_1254_re;
    _T_1255_im <= _T_1254_im;
    _T_1256_re <= _T_1255_re;
    _T_1256_im <= _T_1255_im;
    _T_1257_re <= _T_1256_re;
    _T_1257_im <= _T_1256_im;
    _T_1258_re <= _T_1257_re;
    _T_1258_im <= _T_1257_im;
    _T_1259_re <= _T_1258_re;
    _T_1259_im <= _T_1258_im;
    _T_1260_re <= _T_1259_re;
    _T_1260_im <= _T_1259_im;
    _T_1261_re <= _T_1260_re;
    _T_1261_im <= _T_1260_im;
    _T_1262_re <= _T_1261_re;
    _T_1262_im <= _T_1261_im;
    _T_1263_re <= _T_1262_re;
    _T_1263_im <= _T_1262_im;
    _T_1264_re <= _T_1263_re;
    _T_1264_im <= _T_1263_im;
    _T_1265_re <= _T_1264_re;
    _T_1265_im <= _T_1264_im;
    _T_1266_re <= _T_1265_re;
    _T_1266_im <= _T_1265_im;
    _T_1267_re <= _T_1266_re;
    _T_1267_im <= _T_1266_im;
    _T_1268_re <= _T_1267_re;
    _T_1268_im <= _T_1267_im;
    _T_1269_re <= _T_1268_re;
    _T_1269_im <= _T_1268_im;
    _T_1270_re <= _T_1269_re;
    _T_1270_im <= _T_1269_im;
    _T_1271_re <= _T_1270_re;
    _T_1271_im <= _T_1270_im;
    _T_1272_re <= _T_1271_re;
    _T_1272_im <= _T_1271_im;
    _T_1273_re <= _T_1272_re;
    _T_1273_im <= _T_1272_im;
    _T_1274_re <= _T_1273_re;
    _T_1274_im <= _T_1273_im;
    _T_1275_re <= _T_1274_re;
    _T_1275_im <= _T_1274_im;
    _T_1276_re <= _T_1275_re;
    _T_1276_im <= _T_1275_im;
    _T_1277_re <= _T_1276_re;
    _T_1277_im <= _T_1276_im;
    _T_1278_re <= _T_1277_re;
    _T_1278_im <= _T_1277_im;
    _T_1279_re <= _T_1278_re;
    _T_1279_im <= _T_1278_im;
    _T_1280_re <= _T_1279_re;
    _T_1280_im <= _T_1279_im;
    _T_1281_re <= _T_1280_re;
    _T_1281_im <= _T_1280_im;
    _T_1282_re <= _T_1281_re;
    _T_1282_im <= _T_1281_im;
    _T_1283_re <= _T_1282_re;
    _T_1283_im <= _T_1282_im;
    _T_1284_re <= _T_1283_re;
    _T_1284_im <= _T_1283_im;
    _T_1285_re <= _T_1284_re;
    _T_1285_im <= _T_1284_im;
    _T_1286_re <= _T_1285_re;
    _T_1286_im <= _T_1285_im;
    _T_1287_re <= _T_1286_re;
    _T_1287_im <= _T_1286_im;
    _T_1288_re <= _T_1287_re;
    _T_1288_im <= _T_1287_im;
    _T_1289_re <= _T_1288_re;
    _T_1289_im <= _T_1288_im;
    _T_1290_re <= _T_1289_re;
    _T_1290_im <= _T_1289_im;
    _T_1291_re <= _T_1290_re;
    _T_1291_im <= _T_1290_im;
    _T_1292_re <= _T_1291_re;
    _T_1292_im <= _T_1291_im;
    _T_1293_re <= _T_1292_re;
    _T_1293_im <= _T_1292_im;
    _T_1294_re <= _T_1293_re;
    _T_1294_im <= _T_1293_im;
    _T_1295_re <= _T_1294_re;
    _T_1295_im <= _T_1294_im;
    _T_1296_re <= _T_1295_re;
    _T_1296_im <= _T_1295_im;
    _T_1297_re <= _T_1296_re;
    _T_1297_im <= _T_1296_im;
    _T_1298_re <= _T_1297_re;
    _T_1298_im <= _T_1297_im;
    _T_1299_re <= _T_1298_re;
    _T_1299_im <= _T_1298_im;
    _T_1300_re <= _T_1299_re;
    _T_1300_im <= _T_1299_im;
    _T_1301_re <= _T_1300_re;
    _T_1301_im <= _T_1300_im;
    _T_1302_re <= _T_1301_re;
    _T_1302_im <= _T_1301_im;
    _T_1303_re <= _T_1302_re;
    _T_1303_im <= _T_1302_im;
    _T_1304_re <= _T_1303_re;
    _T_1304_im <= _T_1303_im;
    _T_1305_re <= _T_1304_re;
    _T_1305_im <= _T_1304_im;
    _T_1306_re <= _T_1305_re;
    _T_1306_im <= _T_1305_im;
    _T_1307_re <= _T_1306_re;
    _T_1307_im <= _T_1306_im;
    _T_1308_re <= _T_1307_re;
    _T_1308_im <= _T_1307_im;
    _T_1309_re <= _T_1308_re;
    _T_1309_im <= _T_1308_im;
    _T_1310_re <= _T_1309_re;
    _T_1310_im <= _T_1309_im;
    _T_1311_re <= _T_1310_re;
    _T_1311_im <= _T_1310_im;
    _T_1312_re <= _T_1311_re;
    _T_1312_im <= _T_1311_im;
    _T_1313_re <= _T_1312_re;
    _T_1313_im <= _T_1312_im;
    _T_1314_re <= _T_1313_re;
    _T_1314_im <= _T_1313_im;
    _T_1315_re <= _T_1314_re;
    _T_1315_im <= _T_1314_im;
    _T_1316_re <= _T_1315_re;
    _T_1316_im <= _T_1315_im;
    _T_1317_re <= _T_1316_re;
    _T_1317_im <= _T_1316_im;
    _T_1318_re <= _T_1317_re;
    _T_1318_im <= _T_1317_im;
    _T_1319_re <= _T_1318_re;
    _T_1319_im <= _T_1318_im;
    _T_1320_re <= _T_1319_re;
    _T_1320_im <= _T_1319_im;
    _T_1321_re <= _T_1320_re;
    _T_1321_im <= _T_1320_im;
    _T_1327_re <= Switch_1_io_out1_re;
    _T_1327_im <= Switch_1_io_out1_im;
    _T_1328_re <= _T_1327_re;
    _T_1328_im <= _T_1327_im;
    _T_1329_re <= _T_1328_re;
    _T_1329_im <= _T_1328_im;
    _T_1330_re <= _T_1329_re;
    _T_1330_im <= _T_1329_im;
    _T_1331_re <= _T_1330_re;
    _T_1331_im <= _T_1330_im;
    _T_1332_re <= _T_1331_re;
    _T_1332_im <= _T_1331_im;
    _T_1333_re <= _T_1332_re;
    _T_1333_im <= _T_1332_im;
    _T_1334_re <= _T_1333_re;
    _T_1334_im <= _T_1333_im;
    _T_1335_re <= _T_1334_re;
    _T_1335_im <= _T_1334_im;
    _T_1336_re <= _T_1335_re;
    _T_1336_im <= _T_1335_im;
    _T_1337_re <= _T_1336_re;
    _T_1337_im <= _T_1336_im;
    _T_1338_re <= _T_1337_re;
    _T_1338_im <= _T_1337_im;
    _T_1339_re <= _T_1338_re;
    _T_1339_im <= _T_1338_im;
    _T_1340_re <= _T_1339_re;
    _T_1340_im <= _T_1339_im;
    _T_1341_re <= _T_1340_re;
    _T_1341_im <= _T_1340_im;
    _T_1342_re <= _T_1341_re;
    _T_1342_im <= _T_1341_im;
    _T_1343_re <= _T_1342_re;
    _T_1343_im <= _T_1342_im;
    _T_1344_re <= _T_1343_re;
    _T_1344_im <= _T_1343_im;
    _T_1345_re <= _T_1344_re;
    _T_1345_im <= _T_1344_im;
    _T_1346_re <= _T_1345_re;
    _T_1346_im <= _T_1345_im;
    _T_1347_re <= _T_1346_re;
    _T_1347_im <= _T_1346_im;
    _T_1348_re <= _T_1347_re;
    _T_1348_im <= _T_1347_im;
    _T_1349_re <= _T_1348_re;
    _T_1349_im <= _T_1348_im;
    _T_1350_re <= _T_1349_re;
    _T_1350_im <= _T_1349_im;
    _T_1351_re <= _T_1350_re;
    _T_1351_im <= _T_1350_im;
    _T_1352_re <= _T_1351_re;
    _T_1352_im <= _T_1351_im;
    _T_1353_re <= _T_1352_re;
    _T_1353_im <= _T_1352_im;
    _T_1354_re <= _T_1353_re;
    _T_1354_im <= _T_1353_im;
    _T_1355_re <= _T_1354_re;
    _T_1355_im <= _T_1354_im;
    _T_1356_re <= _T_1355_re;
    _T_1356_im <= _T_1355_im;
    _T_1357_re <= _T_1356_re;
    _T_1357_im <= _T_1356_im;
    _T_1358_re <= _T_1357_re;
    _T_1358_im <= _T_1357_im;
    _T_1359_re <= _T_1358_re;
    _T_1359_im <= _T_1358_im;
    _T_1360_re <= _T_1359_re;
    _T_1360_im <= _T_1359_im;
    _T_1361_re <= _T_1360_re;
    _T_1361_im <= _T_1360_im;
    _T_1362_re <= _T_1361_re;
    _T_1362_im <= _T_1361_im;
    _T_1363_re <= _T_1362_re;
    _T_1363_im <= _T_1362_im;
    _T_1364_re <= _T_1363_re;
    _T_1364_im <= _T_1363_im;
    _T_1365_re <= _T_1364_re;
    _T_1365_im <= _T_1364_im;
    _T_1366_re <= _T_1365_re;
    _T_1366_im <= _T_1365_im;
    _T_1367_re <= _T_1366_re;
    _T_1367_im <= _T_1366_im;
    _T_1368_re <= _T_1367_re;
    _T_1368_im <= _T_1367_im;
    _T_1369_re <= _T_1368_re;
    _T_1369_im <= _T_1368_im;
    _T_1370_re <= _T_1369_re;
    _T_1370_im <= _T_1369_im;
    _T_1371_re <= _T_1370_re;
    _T_1371_im <= _T_1370_im;
    _T_1372_re <= _T_1371_re;
    _T_1372_im <= _T_1371_im;
    _T_1373_re <= _T_1372_re;
    _T_1373_im <= _T_1372_im;
    _T_1374_re <= _T_1373_re;
    _T_1374_im <= _T_1373_im;
    _T_1375_re <= _T_1374_re;
    _T_1375_im <= _T_1374_im;
    _T_1376_re <= _T_1375_re;
    _T_1376_im <= _T_1375_im;
    _T_1377_re <= _T_1376_re;
    _T_1377_im <= _T_1376_im;
    _T_1378_re <= _T_1377_re;
    _T_1378_im <= _T_1377_im;
    _T_1379_re <= _T_1378_re;
    _T_1379_im <= _T_1378_im;
    _T_1380_re <= _T_1379_re;
    _T_1380_im <= _T_1379_im;
    _T_1381_re <= _T_1380_re;
    _T_1381_im <= _T_1380_im;
    _T_1382_re <= _T_1381_re;
    _T_1382_im <= _T_1381_im;
    _T_1383_re <= _T_1382_re;
    _T_1383_im <= _T_1382_im;
    _T_1384_re <= _T_1383_re;
    _T_1384_im <= _T_1383_im;
    _T_1385_re <= _T_1384_re;
    _T_1385_im <= _T_1384_im;
    _T_1386_re <= _T_1385_re;
    _T_1386_im <= _T_1385_im;
    _T_1387_re <= _T_1386_re;
    _T_1387_im <= _T_1386_im;
    _T_1388_re <= _T_1387_re;
    _T_1388_im <= _T_1387_im;
    _T_1389_re <= _T_1388_re;
    _T_1389_im <= _T_1388_im;
    _T_1390_re <= _T_1389_re;
    _T_1390_im <= _T_1389_im;
    _T_1391_re <= _T_1390_re;
    _T_1391_im <= _T_1390_im;
    _T_1392_re <= _T_1391_re;
    _T_1392_im <= _T_1391_im;
    _T_1393_re <= _T_1392_re;
    _T_1393_im <= _T_1392_im;
    _T_1394_re <= _T_1393_re;
    _T_1394_im <= _T_1393_im;
    _T_1395_re <= _T_1394_re;
    _T_1395_im <= _T_1394_im;
    _T_1396_re <= _T_1395_re;
    _T_1396_im <= _T_1395_im;
    _T_1397_re <= _T_1396_re;
    _T_1397_im <= _T_1396_im;
    _T_1398_re <= _T_1397_re;
    _T_1398_im <= _T_1397_im;
    _T_1399_re <= _T_1398_re;
    _T_1399_im <= _T_1398_im;
    _T_1400_re <= _T_1399_re;
    _T_1400_im <= _T_1399_im;
    _T_1401_re <= _T_1400_re;
    _T_1401_im <= _T_1400_im;
    _T_1402_re <= _T_1401_re;
    _T_1402_im <= _T_1401_im;
    _T_1403_re <= _T_1402_re;
    _T_1403_im <= _T_1402_im;
    _T_1404_re <= _T_1403_re;
    _T_1404_im <= _T_1403_im;
    _T_1405_re <= _T_1404_re;
    _T_1405_im <= _T_1404_im;
    _T_1406_re <= _T_1405_re;
    _T_1406_im <= _T_1405_im;
    _T_1407_re <= _T_1406_re;
    _T_1407_im <= _T_1406_im;
    _T_1408_re <= _T_1407_re;
    _T_1408_im <= _T_1407_im;
    _T_1409_re <= _T_1408_re;
    _T_1409_im <= _T_1408_im;
    _T_1410_re <= _T_1409_re;
    _T_1410_im <= _T_1409_im;
    _T_1411_re <= _T_1410_re;
    _T_1411_im <= _T_1410_im;
    _T_1412_re <= _T_1411_re;
    _T_1412_im <= _T_1411_im;
    _T_1413_re <= _T_1412_re;
    _T_1413_im <= _T_1412_im;
    _T_1414_re <= _T_1413_re;
    _T_1414_im <= _T_1413_im;
    _T_1415_re <= _T_1414_re;
    _T_1415_im <= _T_1414_im;
    _T_1416_re <= _T_1415_re;
    _T_1416_im <= _T_1415_im;
    _T_1417_re <= _T_1416_re;
    _T_1417_im <= _T_1416_im;
    _T_1418_re <= _T_1417_re;
    _T_1418_im <= _T_1417_im;
    _T_1419_re <= _T_1418_re;
    _T_1419_im <= _T_1418_im;
    _T_1420_re <= _T_1419_re;
    _T_1420_im <= _T_1419_im;
    _T_1421_re <= _T_1420_re;
    _T_1421_im <= _T_1420_im;
    _T_1422_re <= _T_1421_re;
    _T_1422_im <= _T_1421_im;
    _T_1423_re <= _T_1422_re;
    _T_1423_im <= _T_1422_im;
    _T_1424_re <= _T_1423_re;
    _T_1424_im <= _T_1423_im;
    _T_1425_re <= _T_1424_re;
    _T_1425_im <= _T_1424_im;
    _T_1426_re <= _T_1425_re;
    _T_1426_im <= _T_1425_im;
    _T_1427_re <= _T_1426_re;
    _T_1427_im <= _T_1426_im;
    _T_1428_re <= _T_1427_re;
    _T_1428_im <= _T_1427_im;
    _T_1429_re <= _T_1428_re;
    _T_1429_im <= _T_1428_im;
    _T_1430_re <= _T_1429_re;
    _T_1430_im <= _T_1429_im;
    _T_1431_re <= _T_1430_re;
    _T_1431_im <= _T_1430_im;
    _T_1432_re <= _T_1431_re;
    _T_1432_im <= _T_1431_im;
    _T_1433_re <= _T_1432_re;
    _T_1433_im <= _T_1432_im;
    _T_1434_re <= _T_1433_re;
    _T_1434_im <= _T_1433_im;
    _T_1435_re <= _T_1434_re;
    _T_1435_im <= _T_1434_im;
    _T_1436_re <= _T_1435_re;
    _T_1436_im <= _T_1435_im;
    _T_1437_re <= _T_1436_re;
    _T_1437_im <= _T_1436_im;
    _T_1438_re <= _T_1437_re;
    _T_1438_im <= _T_1437_im;
    _T_1439_re <= _T_1438_re;
    _T_1439_im <= _T_1438_im;
    _T_1440_re <= _T_1439_re;
    _T_1440_im <= _T_1439_im;
    _T_1441_re <= _T_1440_re;
    _T_1441_im <= _T_1440_im;
    _T_1442_re <= _T_1441_re;
    _T_1442_im <= _T_1441_im;
    _T_1443_re <= _T_1442_re;
    _T_1443_im <= _T_1442_im;
    _T_1444_re <= _T_1443_re;
    _T_1444_im <= _T_1443_im;
    _T_1445_re <= _T_1444_re;
    _T_1445_im <= _T_1444_im;
    _T_1446_re <= _T_1445_re;
    _T_1446_im <= _T_1445_im;
    _T_1447_re <= _T_1446_re;
    _T_1447_im <= _T_1446_im;
    _T_1448_re <= _T_1447_re;
    _T_1448_im <= _T_1447_im;
    _T_1449_re <= _T_1448_re;
    _T_1449_im <= _T_1448_im;
    _T_1450_re <= _T_1449_re;
    _T_1450_im <= _T_1449_im;
    _T_1451_re <= _T_1450_re;
    _T_1451_im <= _T_1450_im;
    _T_1452_re <= _T_1451_re;
    _T_1452_im <= _T_1451_im;
    _T_1453_re <= _T_1452_re;
    _T_1453_im <= _T_1452_im;
    _T_1454_re <= _T_1453_re;
    _T_1454_im <= _T_1453_im;
    _T_1457_re <= Butterfly_2_io_out2_re;
    _T_1457_im <= Butterfly_2_io_out2_im;
    _T_1458_re <= _T_1457_re;
    _T_1458_im <= _T_1457_im;
    _T_1459_re <= _T_1458_re;
    _T_1459_im <= _T_1458_im;
    _T_1460_re <= _T_1459_re;
    _T_1460_im <= _T_1459_im;
    _T_1461_re <= _T_1460_re;
    _T_1461_im <= _T_1460_im;
    _T_1462_re <= _T_1461_re;
    _T_1462_im <= _T_1461_im;
    _T_1463_re <= _T_1462_re;
    _T_1463_im <= _T_1462_im;
    _T_1464_re <= _T_1463_re;
    _T_1464_im <= _T_1463_im;
    _T_1465_re <= _T_1464_re;
    _T_1465_im <= _T_1464_im;
    _T_1466_re <= _T_1465_re;
    _T_1466_im <= _T_1465_im;
    _T_1467_re <= _T_1466_re;
    _T_1467_im <= _T_1466_im;
    _T_1468_re <= _T_1467_re;
    _T_1468_im <= _T_1467_im;
    _T_1469_re <= _T_1468_re;
    _T_1469_im <= _T_1468_im;
    _T_1470_re <= _T_1469_re;
    _T_1470_im <= _T_1469_im;
    _T_1471_re <= _T_1470_re;
    _T_1471_im <= _T_1470_im;
    _T_1472_re <= _T_1471_re;
    _T_1472_im <= _T_1471_im;
    _T_1473_re <= _T_1472_re;
    _T_1473_im <= _T_1472_im;
    _T_1474_re <= _T_1473_re;
    _T_1474_im <= _T_1473_im;
    _T_1475_re <= _T_1474_re;
    _T_1475_im <= _T_1474_im;
    _T_1476_re <= _T_1475_re;
    _T_1476_im <= _T_1475_im;
    _T_1477_re <= _T_1476_re;
    _T_1477_im <= _T_1476_im;
    _T_1478_re <= _T_1477_re;
    _T_1478_im <= _T_1477_im;
    _T_1479_re <= _T_1478_re;
    _T_1479_im <= _T_1478_im;
    _T_1480_re <= _T_1479_re;
    _T_1480_im <= _T_1479_im;
    _T_1481_re <= _T_1480_re;
    _T_1481_im <= _T_1480_im;
    _T_1482_re <= _T_1481_re;
    _T_1482_im <= _T_1481_im;
    _T_1483_re <= _T_1482_re;
    _T_1483_im <= _T_1482_im;
    _T_1484_re <= _T_1483_re;
    _T_1484_im <= _T_1483_im;
    _T_1485_re <= _T_1484_re;
    _T_1485_im <= _T_1484_im;
    _T_1486_re <= _T_1485_re;
    _T_1486_im <= _T_1485_im;
    _T_1487_re <= _T_1486_re;
    _T_1487_im <= _T_1486_im;
    _T_1488_re <= _T_1487_re;
    _T_1488_im <= _T_1487_im;
    _T_1489_re <= _T_1488_re;
    _T_1489_im <= _T_1488_im;
    _T_1490_re <= _T_1489_re;
    _T_1490_im <= _T_1489_im;
    _T_1491_re <= _T_1490_re;
    _T_1491_im <= _T_1490_im;
    _T_1492_re <= _T_1491_re;
    _T_1492_im <= _T_1491_im;
    _T_1493_re <= _T_1492_re;
    _T_1493_im <= _T_1492_im;
    _T_1494_re <= _T_1493_re;
    _T_1494_im <= _T_1493_im;
    _T_1495_re <= _T_1494_re;
    _T_1495_im <= _T_1494_im;
    _T_1496_re <= _T_1495_re;
    _T_1496_im <= _T_1495_im;
    _T_1497_re <= _T_1496_re;
    _T_1497_im <= _T_1496_im;
    _T_1498_re <= _T_1497_re;
    _T_1498_im <= _T_1497_im;
    _T_1499_re <= _T_1498_re;
    _T_1499_im <= _T_1498_im;
    _T_1500_re <= _T_1499_re;
    _T_1500_im <= _T_1499_im;
    _T_1501_re <= _T_1500_re;
    _T_1501_im <= _T_1500_im;
    _T_1502_re <= _T_1501_re;
    _T_1502_im <= _T_1501_im;
    _T_1503_re <= _T_1502_re;
    _T_1503_im <= _T_1502_im;
    _T_1504_re <= _T_1503_re;
    _T_1504_im <= _T_1503_im;
    _T_1505_re <= _T_1504_re;
    _T_1505_im <= _T_1504_im;
    _T_1506_re <= _T_1505_re;
    _T_1506_im <= _T_1505_im;
    _T_1507_re <= _T_1506_re;
    _T_1507_im <= _T_1506_im;
    _T_1508_re <= _T_1507_re;
    _T_1508_im <= _T_1507_im;
    _T_1509_re <= _T_1508_re;
    _T_1509_im <= _T_1508_im;
    _T_1510_re <= _T_1509_re;
    _T_1510_im <= _T_1509_im;
    _T_1511_re <= _T_1510_re;
    _T_1511_im <= _T_1510_im;
    _T_1512_re <= _T_1511_re;
    _T_1512_im <= _T_1511_im;
    _T_1513_re <= _T_1512_re;
    _T_1513_im <= _T_1512_im;
    _T_1514_re <= _T_1513_re;
    _T_1514_im <= _T_1513_im;
    _T_1515_re <= _T_1514_re;
    _T_1515_im <= _T_1514_im;
    _T_1516_re <= _T_1515_re;
    _T_1516_im <= _T_1515_im;
    _T_1517_re <= _T_1516_re;
    _T_1517_im <= _T_1516_im;
    _T_1518_re <= _T_1517_re;
    _T_1518_im <= _T_1517_im;
    _T_1519_re <= _T_1518_re;
    _T_1519_im <= _T_1518_im;
    _T_1520_re <= _T_1519_re;
    _T_1520_im <= _T_1519_im;
    _T_1526_re <= Switch_2_io_out1_re;
    _T_1526_im <= Switch_2_io_out1_im;
    _T_1527_re <= _T_1526_re;
    _T_1527_im <= _T_1526_im;
    _T_1528_re <= _T_1527_re;
    _T_1528_im <= _T_1527_im;
    _T_1529_re <= _T_1528_re;
    _T_1529_im <= _T_1528_im;
    _T_1530_re <= _T_1529_re;
    _T_1530_im <= _T_1529_im;
    _T_1531_re <= _T_1530_re;
    _T_1531_im <= _T_1530_im;
    _T_1532_re <= _T_1531_re;
    _T_1532_im <= _T_1531_im;
    _T_1533_re <= _T_1532_re;
    _T_1533_im <= _T_1532_im;
    _T_1534_re <= _T_1533_re;
    _T_1534_im <= _T_1533_im;
    _T_1535_re <= _T_1534_re;
    _T_1535_im <= _T_1534_im;
    _T_1536_re <= _T_1535_re;
    _T_1536_im <= _T_1535_im;
    _T_1537_re <= _T_1536_re;
    _T_1537_im <= _T_1536_im;
    _T_1538_re <= _T_1537_re;
    _T_1538_im <= _T_1537_im;
    _T_1539_re <= _T_1538_re;
    _T_1539_im <= _T_1538_im;
    _T_1540_re <= _T_1539_re;
    _T_1540_im <= _T_1539_im;
    _T_1541_re <= _T_1540_re;
    _T_1541_im <= _T_1540_im;
    _T_1542_re <= _T_1541_re;
    _T_1542_im <= _T_1541_im;
    _T_1543_re <= _T_1542_re;
    _T_1543_im <= _T_1542_im;
    _T_1544_re <= _T_1543_re;
    _T_1544_im <= _T_1543_im;
    _T_1545_re <= _T_1544_re;
    _T_1545_im <= _T_1544_im;
    _T_1546_re <= _T_1545_re;
    _T_1546_im <= _T_1545_im;
    _T_1547_re <= _T_1546_re;
    _T_1547_im <= _T_1546_im;
    _T_1548_re <= _T_1547_re;
    _T_1548_im <= _T_1547_im;
    _T_1549_re <= _T_1548_re;
    _T_1549_im <= _T_1548_im;
    _T_1550_re <= _T_1549_re;
    _T_1550_im <= _T_1549_im;
    _T_1551_re <= _T_1550_re;
    _T_1551_im <= _T_1550_im;
    _T_1552_re <= _T_1551_re;
    _T_1552_im <= _T_1551_im;
    _T_1553_re <= _T_1552_re;
    _T_1553_im <= _T_1552_im;
    _T_1554_re <= _T_1553_re;
    _T_1554_im <= _T_1553_im;
    _T_1555_re <= _T_1554_re;
    _T_1555_im <= _T_1554_im;
    _T_1556_re <= _T_1555_re;
    _T_1556_im <= _T_1555_im;
    _T_1557_re <= _T_1556_re;
    _T_1557_im <= _T_1556_im;
    _T_1558_re <= _T_1557_re;
    _T_1558_im <= _T_1557_im;
    _T_1559_re <= _T_1558_re;
    _T_1559_im <= _T_1558_im;
    _T_1560_re <= _T_1559_re;
    _T_1560_im <= _T_1559_im;
    _T_1561_re <= _T_1560_re;
    _T_1561_im <= _T_1560_im;
    _T_1562_re <= _T_1561_re;
    _T_1562_im <= _T_1561_im;
    _T_1563_re <= _T_1562_re;
    _T_1563_im <= _T_1562_im;
    _T_1564_re <= _T_1563_re;
    _T_1564_im <= _T_1563_im;
    _T_1565_re <= _T_1564_re;
    _T_1565_im <= _T_1564_im;
    _T_1566_re <= _T_1565_re;
    _T_1566_im <= _T_1565_im;
    _T_1567_re <= _T_1566_re;
    _T_1567_im <= _T_1566_im;
    _T_1568_re <= _T_1567_re;
    _T_1568_im <= _T_1567_im;
    _T_1569_re <= _T_1568_re;
    _T_1569_im <= _T_1568_im;
    _T_1570_re <= _T_1569_re;
    _T_1570_im <= _T_1569_im;
    _T_1571_re <= _T_1570_re;
    _T_1571_im <= _T_1570_im;
    _T_1572_re <= _T_1571_re;
    _T_1572_im <= _T_1571_im;
    _T_1573_re <= _T_1572_re;
    _T_1573_im <= _T_1572_im;
    _T_1574_re <= _T_1573_re;
    _T_1574_im <= _T_1573_im;
    _T_1575_re <= _T_1574_re;
    _T_1575_im <= _T_1574_im;
    _T_1576_re <= _T_1575_re;
    _T_1576_im <= _T_1575_im;
    _T_1577_re <= _T_1576_re;
    _T_1577_im <= _T_1576_im;
    _T_1578_re <= _T_1577_re;
    _T_1578_im <= _T_1577_im;
    _T_1579_re <= _T_1578_re;
    _T_1579_im <= _T_1578_im;
    _T_1580_re <= _T_1579_re;
    _T_1580_im <= _T_1579_im;
    _T_1581_re <= _T_1580_re;
    _T_1581_im <= _T_1580_im;
    _T_1582_re <= _T_1581_re;
    _T_1582_im <= _T_1581_im;
    _T_1583_re <= _T_1582_re;
    _T_1583_im <= _T_1582_im;
    _T_1584_re <= _T_1583_re;
    _T_1584_im <= _T_1583_im;
    _T_1585_re <= _T_1584_re;
    _T_1585_im <= _T_1584_im;
    _T_1586_re <= _T_1585_re;
    _T_1586_im <= _T_1585_im;
    _T_1587_re <= _T_1586_re;
    _T_1587_im <= _T_1586_im;
    _T_1588_re <= _T_1587_re;
    _T_1588_im <= _T_1587_im;
    _T_1589_re <= _T_1588_re;
    _T_1589_im <= _T_1588_im;
    _T_1592_re <= Butterfly_3_io_out2_re;
    _T_1592_im <= Butterfly_3_io_out2_im;
    _T_1593_re <= _T_1592_re;
    _T_1593_im <= _T_1592_im;
    _T_1594_re <= _T_1593_re;
    _T_1594_im <= _T_1593_im;
    _T_1595_re <= _T_1594_re;
    _T_1595_im <= _T_1594_im;
    _T_1596_re <= _T_1595_re;
    _T_1596_im <= _T_1595_im;
    _T_1597_re <= _T_1596_re;
    _T_1597_im <= _T_1596_im;
    _T_1598_re <= _T_1597_re;
    _T_1598_im <= _T_1597_im;
    _T_1599_re <= _T_1598_re;
    _T_1599_im <= _T_1598_im;
    _T_1600_re <= _T_1599_re;
    _T_1600_im <= _T_1599_im;
    _T_1601_re <= _T_1600_re;
    _T_1601_im <= _T_1600_im;
    _T_1602_re <= _T_1601_re;
    _T_1602_im <= _T_1601_im;
    _T_1603_re <= _T_1602_re;
    _T_1603_im <= _T_1602_im;
    _T_1604_re <= _T_1603_re;
    _T_1604_im <= _T_1603_im;
    _T_1605_re <= _T_1604_re;
    _T_1605_im <= _T_1604_im;
    _T_1606_re <= _T_1605_re;
    _T_1606_im <= _T_1605_im;
    _T_1607_re <= _T_1606_re;
    _T_1607_im <= _T_1606_im;
    _T_1608_re <= _T_1607_re;
    _T_1608_im <= _T_1607_im;
    _T_1609_re <= _T_1608_re;
    _T_1609_im <= _T_1608_im;
    _T_1610_re <= _T_1609_re;
    _T_1610_im <= _T_1609_im;
    _T_1611_re <= _T_1610_re;
    _T_1611_im <= _T_1610_im;
    _T_1612_re <= _T_1611_re;
    _T_1612_im <= _T_1611_im;
    _T_1613_re <= _T_1612_re;
    _T_1613_im <= _T_1612_im;
    _T_1614_re <= _T_1613_re;
    _T_1614_im <= _T_1613_im;
    _T_1615_re <= _T_1614_re;
    _T_1615_im <= _T_1614_im;
    _T_1616_re <= _T_1615_re;
    _T_1616_im <= _T_1615_im;
    _T_1617_re <= _T_1616_re;
    _T_1617_im <= _T_1616_im;
    _T_1618_re <= _T_1617_re;
    _T_1618_im <= _T_1617_im;
    _T_1619_re <= _T_1618_re;
    _T_1619_im <= _T_1618_im;
    _T_1620_re <= _T_1619_re;
    _T_1620_im <= _T_1619_im;
    _T_1621_re <= _T_1620_re;
    _T_1621_im <= _T_1620_im;
    _T_1622_re <= _T_1621_re;
    _T_1622_im <= _T_1621_im;
    _T_1623_re <= _T_1622_re;
    _T_1623_im <= _T_1622_im;
    _T_1629_re <= Switch_3_io_out1_re;
    _T_1629_im <= Switch_3_io_out1_im;
    _T_1630_re <= _T_1629_re;
    _T_1630_im <= _T_1629_im;
    _T_1631_re <= _T_1630_re;
    _T_1631_im <= _T_1630_im;
    _T_1632_re <= _T_1631_re;
    _T_1632_im <= _T_1631_im;
    _T_1633_re <= _T_1632_re;
    _T_1633_im <= _T_1632_im;
    _T_1634_re <= _T_1633_re;
    _T_1634_im <= _T_1633_im;
    _T_1635_re <= _T_1634_re;
    _T_1635_im <= _T_1634_im;
    _T_1636_re <= _T_1635_re;
    _T_1636_im <= _T_1635_im;
    _T_1637_re <= _T_1636_re;
    _T_1637_im <= _T_1636_im;
    _T_1638_re <= _T_1637_re;
    _T_1638_im <= _T_1637_im;
    _T_1639_re <= _T_1638_re;
    _T_1639_im <= _T_1638_im;
    _T_1640_re <= _T_1639_re;
    _T_1640_im <= _T_1639_im;
    _T_1641_re <= _T_1640_re;
    _T_1641_im <= _T_1640_im;
    _T_1642_re <= _T_1641_re;
    _T_1642_im <= _T_1641_im;
    _T_1643_re <= _T_1642_re;
    _T_1643_im <= _T_1642_im;
    _T_1644_re <= _T_1643_re;
    _T_1644_im <= _T_1643_im;
    _T_1645_re <= _T_1644_re;
    _T_1645_im <= _T_1644_im;
    _T_1646_re <= _T_1645_re;
    _T_1646_im <= _T_1645_im;
    _T_1647_re <= _T_1646_re;
    _T_1647_im <= _T_1646_im;
    _T_1648_re <= _T_1647_re;
    _T_1648_im <= _T_1647_im;
    _T_1649_re <= _T_1648_re;
    _T_1649_im <= _T_1648_im;
    _T_1650_re <= _T_1649_re;
    _T_1650_im <= _T_1649_im;
    _T_1651_re <= _T_1650_re;
    _T_1651_im <= _T_1650_im;
    _T_1652_re <= _T_1651_re;
    _T_1652_im <= _T_1651_im;
    _T_1653_re <= _T_1652_re;
    _T_1653_im <= _T_1652_im;
    _T_1654_re <= _T_1653_re;
    _T_1654_im <= _T_1653_im;
    _T_1655_re <= _T_1654_re;
    _T_1655_im <= _T_1654_im;
    _T_1656_re <= _T_1655_re;
    _T_1656_im <= _T_1655_im;
    _T_1657_re <= _T_1656_re;
    _T_1657_im <= _T_1656_im;
    _T_1658_re <= _T_1657_re;
    _T_1658_im <= _T_1657_im;
    _T_1659_re <= _T_1658_re;
    _T_1659_im <= _T_1658_im;
    _T_1660_re <= _T_1659_re;
    _T_1660_im <= _T_1659_im;
    _T_1663_re <= Butterfly_4_io_out2_re;
    _T_1663_im <= Butterfly_4_io_out2_im;
    _T_1664_re <= _T_1663_re;
    _T_1664_im <= _T_1663_im;
    _T_1665_re <= _T_1664_re;
    _T_1665_im <= _T_1664_im;
    _T_1666_re <= _T_1665_re;
    _T_1666_im <= _T_1665_im;
    _T_1667_re <= _T_1666_re;
    _T_1667_im <= _T_1666_im;
    _T_1668_re <= _T_1667_re;
    _T_1668_im <= _T_1667_im;
    _T_1669_re <= _T_1668_re;
    _T_1669_im <= _T_1668_im;
    _T_1670_re <= _T_1669_re;
    _T_1670_im <= _T_1669_im;
    _T_1671_re <= _T_1670_re;
    _T_1671_im <= _T_1670_im;
    _T_1672_re <= _T_1671_re;
    _T_1672_im <= _T_1671_im;
    _T_1673_re <= _T_1672_re;
    _T_1673_im <= _T_1672_im;
    _T_1674_re <= _T_1673_re;
    _T_1674_im <= _T_1673_im;
    _T_1675_re <= _T_1674_re;
    _T_1675_im <= _T_1674_im;
    _T_1676_re <= _T_1675_re;
    _T_1676_im <= _T_1675_im;
    _T_1677_re <= _T_1676_re;
    _T_1677_im <= _T_1676_im;
    _T_1678_re <= _T_1677_re;
    _T_1678_im <= _T_1677_im;
    _T_1684_re <= Switch_4_io_out1_re;
    _T_1684_im <= Switch_4_io_out1_im;
    _T_1685_re <= _T_1684_re;
    _T_1685_im <= _T_1684_im;
    _T_1686_re <= _T_1685_re;
    _T_1686_im <= _T_1685_im;
    _T_1687_re <= _T_1686_re;
    _T_1687_im <= _T_1686_im;
    _T_1688_re <= _T_1687_re;
    _T_1688_im <= _T_1687_im;
    _T_1689_re <= _T_1688_re;
    _T_1689_im <= _T_1688_im;
    _T_1690_re <= _T_1689_re;
    _T_1690_im <= _T_1689_im;
    _T_1691_re <= _T_1690_re;
    _T_1691_im <= _T_1690_im;
    _T_1692_re <= _T_1691_re;
    _T_1692_im <= _T_1691_im;
    _T_1693_re <= _T_1692_re;
    _T_1693_im <= _T_1692_im;
    _T_1694_re <= _T_1693_re;
    _T_1694_im <= _T_1693_im;
    _T_1695_re <= _T_1694_re;
    _T_1695_im <= _T_1694_im;
    _T_1696_re <= _T_1695_re;
    _T_1696_im <= _T_1695_im;
    _T_1697_re <= _T_1696_re;
    _T_1697_im <= _T_1696_im;
    _T_1698_re <= _T_1697_re;
    _T_1698_im <= _T_1697_im;
    _T_1699_re <= _T_1698_re;
    _T_1699_im <= _T_1698_im;
    _T_1702_re <= Butterfly_5_io_out2_re;
    _T_1702_im <= Butterfly_5_io_out2_im;
    _T_1703_re <= _T_1702_re;
    _T_1703_im <= _T_1702_im;
    _T_1704_re <= _T_1703_re;
    _T_1704_im <= _T_1703_im;
    _T_1705_re <= _T_1704_re;
    _T_1705_im <= _T_1704_im;
    _T_1706_re <= _T_1705_re;
    _T_1706_im <= _T_1705_im;
    _T_1707_re <= _T_1706_re;
    _T_1707_im <= _T_1706_im;
    _T_1708_re <= _T_1707_re;
    _T_1708_im <= _T_1707_im;
    _T_1709_re <= _T_1708_re;
    _T_1709_im <= _T_1708_im;
    _T_1715_re <= Switch_5_io_out1_re;
    _T_1715_im <= Switch_5_io_out1_im;
    _T_1716_re <= _T_1715_re;
    _T_1716_im <= _T_1715_im;
    _T_1717_re <= _T_1716_re;
    _T_1717_im <= _T_1716_im;
    _T_1718_re <= _T_1717_re;
    _T_1718_im <= _T_1717_im;
    _T_1719_re <= _T_1718_re;
    _T_1719_im <= _T_1718_im;
    _T_1720_re <= _T_1719_re;
    _T_1720_im <= _T_1719_im;
    _T_1721_re <= _T_1720_re;
    _T_1721_im <= _T_1720_im;
    _T_1722_re <= _T_1721_re;
    _T_1722_im <= _T_1721_im;
    _T_1725_re <= Butterfly_6_io_out2_re;
    _T_1725_im <= Butterfly_6_io_out2_im;
    _T_1726_re <= _T_1725_re;
    _T_1726_im <= _T_1725_im;
    _T_1727_re <= _T_1726_re;
    _T_1727_im <= _T_1726_im;
    _T_1728_re <= _T_1727_re;
    _T_1728_im <= _T_1727_im;
    _T_1734_re <= Switch_6_io_out1_re;
    _T_1734_im <= Switch_6_io_out1_im;
    _T_1735_re <= _T_1734_re;
    _T_1735_im <= _T_1734_im;
    _T_1736_re <= _T_1735_re;
    _T_1736_im <= _T_1735_im;
    _T_1737_re <= _T_1736_re;
    _T_1737_im <= _T_1736_im;
    _T_1740_re <= Butterfly_7_io_out2_re;
    _T_1740_im <= Butterfly_7_io_out2_im;
    _T_1741_re <= _T_1740_re;
    _T_1741_im <= _T_1740_im;
    _T_1747_re <= Switch_7_io_out1_re;
    _T_1747_im <= Switch_7_io_out1_im;
    _T_1748_re <= _T_1747_re;
    _T_1748_im <= _T_1747_im;
    _T_1751_re <= Butterfly_8_io_out2_re;
    _T_1751_im <= Butterfly_8_io_out2_im;
    out1D1_re <= Switch_8_io_out1_re;
    out1D1_im <= Switch_8_io_out1_im;
    _T_1752_re <= ComplexAdd_io_res_re;
    _T_1752_im <= ComplexAdd_io_res_im;
    _T_1753_re <= ComplexSub_io_res_re;
    _T_1753_im <= ComplexSub_io_res_im;
  end
endmodule
