module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T; // @[Butterfly.scala 57:28]
  wire [63:0] _T_1; // @[Butterfly.scala 57:52]
  wire [63:0] _T_4; // @[Butterfly.scala 57:40]
  wire [63:0] _T_5; // @[Butterfly.scala 58:28]
  wire [63:0] _T_6; // @[Butterfly.scala 58:52]
  wire [63:0] _T_9; // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2; // @[Butterfly.scala 58:15]
  assign _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  assign _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  assign _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  assign _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  assign _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  assign _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  assign _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT256(
    input clk_in1_p,
    input clk_in1_n,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
    wire clock;
    clk_wiz_0 clk_wiz_0_inst0
       (
        // Clock out ports
        .clk_out1(clock),     // output clk_out1
       // Clock in ports
        .clk_in1_p(clk_in1_p),    // input clk_in1_p
        .clk_in1_n(clk_in1_n));    // input clk_in1_n
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [7:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [7:0] _T_1; // @[FFT.scala 42:16]
  wire [31:0] _GEN_2; // @[FFT.scala 34:12]
  wire [31:0] _GEN_3; // @[FFT.scala 34:12]
  wire [31:0] _GEN_4; // @[FFT.scala 34:12]
  wire [31:0] _GEN_5; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6; // @[FFT.scala 34:12]
  wire [31:0] _GEN_7; // @[FFT.scala 34:12]
  wire [31:0] _GEN_8; // @[FFT.scala 34:12]
  wire [31:0] _GEN_9; // @[FFT.scala 34:12]
  wire [31:0] _GEN_10; // @[FFT.scala 34:12]
  wire [31:0] _GEN_11; // @[FFT.scala 34:12]
  wire [31:0] _GEN_12; // @[FFT.scala 34:12]
  wire [31:0] _GEN_13; // @[FFT.scala 34:12]
  wire [31:0] _GEN_14; // @[FFT.scala 34:12]
  wire [31:0] _GEN_15; // @[FFT.scala 34:12]
  wire [31:0] _GEN_16; // @[FFT.scala 34:12]
  wire [31:0] _GEN_17; // @[FFT.scala 34:12]
  wire [31:0] _GEN_18; // @[FFT.scala 34:12]
  wire [31:0] _GEN_19; // @[FFT.scala 34:12]
  wire [31:0] _GEN_20; // @[FFT.scala 34:12]
  wire [31:0] _GEN_21; // @[FFT.scala 34:12]
  wire [31:0] _GEN_22; // @[FFT.scala 34:12]
  wire [31:0] _GEN_23; // @[FFT.scala 34:12]
  wire [31:0] _GEN_24; // @[FFT.scala 34:12]
  wire [31:0] _GEN_25; // @[FFT.scala 34:12]
  wire [31:0] _GEN_26; // @[FFT.scala 34:12]
  wire [31:0] _GEN_27; // @[FFT.scala 34:12]
  wire [31:0] _GEN_28; // @[FFT.scala 34:12]
  wire [31:0] _GEN_29; // @[FFT.scala 34:12]
  wire [31:0] _GEN_30; // @[FFT.scala 34:12]
  wire [31:0] _GEN_31; // @[FFT.scala 34:12]
  wire [31:0] _GEN_32; // @[FFT.scala 34:12]
  wire [31:0] _GEN_33; // @[FFT.scala 34:12]
  wire [31:0] _GEN_34; // @[FFT.scala 34:12]
  wire [31:0] _GEN_35; // @[FFT.scala 34:12]
  wire [31:0] _GEN_36; // @[FFT.scala 34:12]
  wire [31:0] _GEN_37; // @[FFT.scala 34:12]
  wire [31:0] _GEN_38; // @[FFT.scala 34:12]
  wire [31:0] _GEN_39; // @[FFT.scala 34:12]
  wire [31:0] _GEN_40; // @[FFT.scala 34:12]
  wire [31:0] _GEN_41; // @[FFT.scala 34:12]
  wire [31:0] _GEN_42; // @[FFT.scala 34:12]
  wire [31:0] _GEN_43; // @[FFT.scala 34:12]
  wire [31:0] _GEN_44; // @[FFT.scala 34:12]
  wire [31:0] _GEN_45; // @[FFT.scala 34:12]
  wire [31:0] _GEN_46; // @[FFT.scala 34:12]
  wire [31:0] _GEN_47; // @[FFT.scala 34:12]
  wire [31:0] _GEN_48; // @[FFT.scala 34:12]
  wire [31:0] _GEN_49; // @[FFT.scala 34:12]
  wire [31:0] _GEN_50; // @[FFT.scala 34:12]
  wire [31:0] _GEN_51; // @[FFT.scala 34:12]
  wire [31:0] _GEN_52; // @[FFT.scala 34:12]
  wire [31:0] _GEN_53; // @[FFT.scala 34:12]
  wire [31:0] _GEN_54; // @[FFT.scala 34:12]
  wire [31:0] _GEN_55; // @[FFT.scala 34:12]
  wire [31:0] _GEN_56; // @[FFT.scala 34:12]
  wire [31:0] _GEN_57; // @[FFT.scala 34:12]
  wire [31:0] _GEN_58; // @[FFT.scala 34:12]
  wire [31:0] _GEN_59; // @[FFT.scala 34:12]
  wire [31:0] _GEN_60; // @[FFT.scala 34:12]
  wire [31:0] _GEN_61; // @[FFT.scala 34:12]
  wire [31:0] _GEN_62; // @[FFT.scala 34:12]
  wire [31:0] _GEN_63; // @[FFT.scala 34:12]
  wire [31:0] _GEN_64; // @[FFT.scala 34:12]
  wire [31:0] _GEN_65; // @[FFT.scala 34:12]
  wire [31:0] _GEN_66; // @[FFT.scala 34:12]
  wire [31:0] _GEN_67; // @[FFT.scala 34:12]
  wire [31:0] _GEN_68; // @[FFT.scala 34:12]
  wire [31:0] _GEN_69; // @[FFT.scala 34:12]
  wire [31:0] _GEN_70; // @[FFT.scala 34:12]
  wire [31:0] _GEN_71; // @[FFT.scala 34:12]
  wire [31:0] _GEN_72; // @[FFT.scala 34:12]
  wire [31:0] _GEN_73; // @[FFT.scala 34:12]
  wire [31:0] _GEN_74; // @[FFT.scala 34:12]
  wire [31:0] _GEN_75; // @[FFT.scala 34:12]
  wire [31:0] _GEN_76; // @[FFT.scala 34:12]
  wire [31:0] _GEN_77; // @[FFT.scala 34:12]
  wire [31:0] _GEN_78; // @[FFT.scala 34:12]
  wire [31:0] _GEN_79; // @[FFT.scala 34:12]
  wire [31:0] _GEN_80; // @[FFT.scala 34:12]
  wire [31:0] _GEN_81; // @[FFT.scala 34:12]
  wire [31:0] _GEN_82; // @[FFT.scala 34:12]
  wire [31:0] _GEN_83; // @[FFT.scala 34:12]
  wire [31:0] _GEN_84; // @[FFT.scala 34:12]
  wire [31:0] _GEN_85; // @[FFT.scala 34:12]
  wire [31:0] _GEN_86; // @[FFT.scala 34:12]
  wire [31:0] _GEN_87; // @[FFT.scala 34:12]
  wire [31:0] _GEN_88; // @[FFT.scala 34:12]
  wire [31:0] _GEN_89; // @[FFT.scala 34:12]
  wire [31:0] _GEN_90; // @[FFT.scala 34:12]
  wire [31:0] _GEN_91; // @[FFT.scala 34:12]
  wire [31:0] _GEN_92; // @[FFT.scala 34:12]
  wire [31:0] _GEN_93; // @[FFT.scala 34:12]
  wire [31:0] _GEN_94; // @[FFT.scala 34:12]
  wire [31:0] _GEN_95; // @[FFT.scala 34:12]
  wire [31:0] _GEN_96; // @[FFT.scala 34:12]
  wire [31:0] _GEN_97; // @[FFT.scala 34:12]
  wire [31:0] _GEN_98; // @[FFT.scala 34:12]
  wire [31:0] _GEN_99; // @[FFT.scala 34:12]
  wire [31:0] _GEN_100; // @[FFT.scala 34:12]
  wire [31:0] _GEN_101; // @[FFT.scala 34:12]
  wire [31:0] _GEN_102; // @[FFT.scala 34:12]
  wire [31:0] _GEN_103; // @[FFT.scala 34:12]
  wire [31:0] _GEN_104; // @[FFT.scala 34:12]
  wire [31:0] _GEN_105; // @[FFT.scala 34:12]
  wire [31:0] _GEN_106; // @[FFT.scala 34:12]
  wire [31:0] _GEN_107; // @[FFT.scala 34:12]
  wire [31:0] _GEN_108; // @[FFT.scala 34:12]
  wire [31:0] _GEN_109; // @[FFT.scala 34:12]
  wire [31:0] _GEN_110; // @[FFT.scala 34:12]
  wire [31:0] _GEN_111; // @[FFT.scala 34:12]
  wire [31:0] _GEN_112; // @[FFT.scala 34:12]
  wire [31:0] _GEN_113; // @[FFT.scala 34:12]
  wire [31:0] _GEN_114; // @[FFT.scala 34:12]
  wire [31:0] _GEN_115; // @[FFT.scala 34:12]
  wire [31:0] _GEN_116; // @[FFT.scala 34:12]
  wire [31:0] _GEN_117; // @[FFT.scala 34:12]
  wire [31:0] _GEN_118; // @[FFT.scala 34:12]
  wire [31:0] _GEN_119; // @[FFT.scala 34:12]
  wire [31:0] _GEN_120; // @[FFT.scala 34:12]
  wire [31:0] _GEN_121; // @[FFT.scala 34:12]
  wire [31:0] _GEN_122; // @[FFT.scala 34:12]
  wire [31:0] _GEN_123; // @[FFT.scala 34:12]
  wire [31:0] _GEN_124; // @[FFT.scala 34:12]
  wire [31:0] _GEN_125; // @[FFT.scala 34:12]
  wire [31:0] _GEN_126; // @[FFT.scala 34:12]
  wire [31:0] _GEN_127; // @[FFT.scala 34:12]
  wire [31:0] _GEN_130; // @[FFT.scala 35:12]
  wire [31:0] _GEN_131; // @[FFT.scala 35:12]
  wire [31:0] _GEN_132; // @[FFT.scala 35:12]
  wire [31:0] _GEN_133; // @[FFT.scala 35:12]
  wire [31:0] _GEN_134; // @[FFT.scala 35:12]
  wire [31:0] _GEN_135; // @[FFT.scala 35:12]
  wire [31:0] _GEN_136; // @[FFT.scala 35:12]
  wire [31:0] _GEN_137; // @[FFT.scala 35:12]
  wire [31:0] _GEN_138; // @[FFT.scala 35:12]
  wire [31:0] _GEN_139; // @[FFT.scala 35:12]
  wire [31:0] _GEN_140; // @[FFT.scala 35:12]
  wire [31:0] _GEN_141; // @[FFT.scala 35:12]
  wire [31:0] _GEN_142; // @[FFT.scala 35:12]
  wire [31:0] _GEN_143; // @[FFT.scala 35:12]
  wire [31:0] _GEN_144; // @[FFT.scala 35:12]
  wire [31:0] _GEN_145; // @[FFT.scala 35:12]
  wire [31:0] _GEN_146; // @[FFT.scala 35:12]
  wire [31:0] _GEN_147; // @[FFT.scala 35:12]
  wire [31:0] _GEN_148; // @[FFT.scala 35:12]
  wire [31:0] _GEN_149; // @[FFT.scala 35:12]
  wire [31:0] _GEN_150; // @[FFT.scala 35:12]
  wire [31:0] _GEN_151; // @[FFT.scala 35:12]
  wire [31:0] _GEN_152; // @[FFT.scala 35:12]
  wire [31:0] _GEN_153; // @[FFT.scala 35:12]
  wire [31:0] _GEN_154; // @[FFT.scala 35:12]
  wire [31:0] _GEN_155; // @[FFT.scala 35:12]
  wire [31:0] _GEN_156; // @[FFT.scala 35:12]
  wire [31:0] _GEN_157; // @[FFT.scala 35:12]
  wire [31:0] _GEN_158; // @[FFT.scala 35:12]
  wire [31:0] _GEN_159; // @[FFT.scala 35:12]
  wire [31:0] _GEN_160; // @[FFT.scala 35:12]
  wire [31:0] _GEN_161; // @[FFT.scala 35:12]
  wire [31:0] _GEN_162; // @[FFT.scala 35:12]
  wire [31:0] _GEN_163; // @[FFT.scala 35:12]
  wire [31:0] _GEN_164; // @[FFT.scala 35:12]
  wire [31:0] _GEN_165; // @[FFT.scala 35:12]
  wire [31:0] _GEN_166; // @[FFT.scala 35:12]
  wire [31:0] _GEN_167; // @[FFT.scala 35:12]
  wire [31:0] _GEN_168; // @[FFT.scala 35:12]
  wire [31:0] _GEN_169; // @[FFT.scala 35:12]
  wire [31:0] _GEN_170; // @[FFT.scala 35:12]
  wire [31:0] _GEN_171; // @[FFT.scala 35:12]
  wire [31:0] _GEN_172; // @[FFT.scala 35:12]
  wire [31:0] _GEN_173; // @[FFT.scala 35:12]
  wire [31:0] _GEN_174; // @[FFT.scala 35:12]
  wire [31:0] _GEN_175; // @[FFT.scala 35:12]
  wire [31:0] _GEN_176; // @[FFT.scala 35:12]
  wire [31:0] _GEN_177; // @[FFT.scala 35:12]
  wire [31:0] _GEN_178; // @[FFT.scala 35:12]
  wire [31:0] _GEN_179; // @[FFT.scala 35:12]
  wire [31:0] _GEN_180; // @[FFT.scala 35:12]
  wire [31:0] _GEN_181; // @[FFT.scala 35:12]
  wire [31:0] _GEN_182; // @[FFT.scala 35:12]
  wire [31:0] _GEN_183; // @[FFT.scala 35:12]
  wire [31:0] _GEN_184; // @[FFT.scala 35:12]
  wire [31:0] _GEN_185; // @[FFT.scala 35:12]
  wire [31:0] _GEN_186; // @[FFT.scala 35:12]
  wire [31:0] _GEN_187; // @[FFT.scala 35:12]
  wire [31:0] _GEN_188; // @[FFT.scala 35:12]
  wire [31:0] _GEN_189; // @[FFT.scala 35:12]
  wire [31:0] _GEN_190; // @[FFT.scala 35:12]
  wire [31:0] _GEN_191; // @[FFT.scala 35:12]
  wire [31:0] _GEN_192; // @[FFT.scala 35:12]
  wire [31:0] _GEN_193; // @[FFT.scala 35:12]
  wire [31:0] _GEN_194; // @[FFT.scala 35:12]
  wire [31:0] _GEN_195; // @[FFT.scala 35:12]
  wire [31:0] _GEN_196; // @[FFT.scala 35:12]
  wire [31:0] _GEN_197; // @[FFT.scala 35:12]
  wire [31:0] _GEN_198; // @[FFT.scala 35:12]
  wire [31:0] _GEN_199; // @[FFT.scala 35:12]
  wire [31:0] _GEN_200; // @[FFT.scala 35:12]
  wire [31:0] _GEN_201; // @[FFT.scala 35:12]
  wire [31:0] _GEN_202; // @[FFT.scala 35:12]
  wire [31:0] _GEN_203; // @[FFT.scala 35:12]
  wire [31:0] _GEN_204; // @[FFT.scala 35:12]
  wire [31:0] _GEN_205; // @[FFT.scala 35:12]
  wire [31:0] _GEN_206; // @[FFT.scala 35:12]
  wire [31:0] _GEN_207; // @[FFT.scala 35:12]
  wire [31:0] _GEN_208; // @[FFT.scala 35:12]
  wire [31:0] _GEN_209; // @[FFT.scala 35:12]
  wire [31:0] _GEN_210; // @[FFT.scala 35:12]
  wire [31:0] _GEN_211; // @[FFT.scala 35:12]
  wire [31:0] _GEN_212; // @[FFT.scala 35:12]
  wire [31:0] _GEN_213; // @[FFT.scala 35:12]
  wire [31:0] _GEN_214; // @[FFT.scala 35:12]
  wire [31:0] _GEN_215; // @[FFT.scala 35:12]
  wire [31:0] _GEN_216; // @[FFT.scala 35:12]
  wire [31:0] _GEN_217; // @[FFT.scala 35:12]
  wire [31:0] _GEN_218; // @[FFT.scala 35:12]
  wire [31:0] _GEN_219; // @[FFT.scala 35:12]
  wire [31:0] _GEN_220; // @[FFT.scala 35:12]
  wire [31:0] _GEN_221; // @[FFT.scala 35:12]
  wire [31:0] _GEN_222; // @[FFT.scala 35:12]
  wire [31:0] _GEN_223; // @[FFT.scala 35:12]
  wire [31:0] _GEN_224; // @[FFT.scala 35:12]
  wire [31:0] _GEN_225; // @[FFT.scala 35:12]
  wire [31:0] _GEN_226; // @[FFT.scala 35:12]
  wire [31:0] _GEN_227; // @[FFT.scala 35:12]
  wire [31:0] _GEN_228; // @[FFT.scala 35:12]
  wire [31:0] _GEN_229; // @[FFT.scala 35:12]
  wire [31:0] _GEN_230; // @[FFT.scala 35:12]
  wire [31:0] _GEN_231; // @[FFT.scala 35:12]
  wire [31:0] _GEN_232; // @[FFT.scala 35:12]
  wire [31:0] _GEN_233; // @[FFT.scala 35:12]
  wire [31:0] _GEN_234; // @[FFT.scala 35:12]
  wire [31:0] _GEN_235; // @[FFT.scala 35:12]
  wire [31:0] _GEN_236; // @[FFT.scala 35:12]
  wire [31:0] _GEN_237; // @[FFT.scala 35:12]
  wire [31:0] _GEN_238; // @[FFT.scala 35:12]
  wire [31:0] _GEN_239; // @[FFT.scala 35:12]
  wire [31:0] _GEN_240; // @[FFT.scala 35:12]
  wire [31:0] _GEN_241; // @[FFT.scala 35:12]
  wire [31:0] _GEN_242; // @[FFT.scala 35:12]
  wire [31:0] _GEN_243; // @[FFT.scala 35:12]
  wire [31:0] _GEN_244; // @[FFT.scala 35:12]
  wire [31:0] _GEN_245; // @[FFT.scala 35:12]
  wire [31:0] _GEN_246; // @[FFT.scala 35:12]
  wire [31:0] _GEN_247; // @[FFT.scala 35:12]
  wire [31:0] _GEN_248; // @[FFT.scala 35:12]
  wire [31:0] _GEN_249; // @[FFT.scala 35:12]
  wire [31:0] _GEN_250; // @[FFT.scala 35:12]
  wire [31:0] _GEN_251; // @[FFT.scala 35:12]
  wire [31:0] _GEN_252; // @[FFT.scala 35:12]
  wire [31:0] _GEN_253; // @[FFT.scala 35:12]
  wire [31:0] _GEN_254; // @[FFT.scala 35:12]
  wire [31:0] _GEN_255; // @[FFT.scala 35:12]
  reg [31:0] _T_132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [31:0] _T_132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [31:0] _T_133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [31:0] _T_133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] _T_134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [31:0] _T_134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [31:0] _T_135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  wire [31:0] _GEN_642; // @[FFT.scala 34:12]
  wire [31:0] _GEN_643; // @[FFT.scala 34:12]
  wire [31:0] _GEN_644; // @[FFT.scala 34:12]
  wire [31:0] _GEN_645; // @[FFT.scala 34:12]
  wire [31:0] _GEN_646; // @[FFT.scala 34:12]
  wire [31:0] _GEN_647; // @[FFT.scala 34:12]
  wire [31:0] _GEN_648; // @[FFT.scala 34:12]
  wire [31:0] _GEN_649; // @[FFT.scala 34:12]
  wire [31:0] _GEN_650; // @[FFT.scala 34:12]
  wire [31:0] _GEN_651; // @[FFT.scala 34:12]
  wire [31:0] _GEN_652; // @[FFT.scala 34:12]
  wire [31:0] _GEN_653; // @[FFT.scala 34:12]
  wire [31:0] _GEN_654; // @[FFT.scala 34:12]
  wire [31:0] _GEN_655; // @[FFT.scala 34:12]
  wire [31:0] _GEN_656; // @[FFT.scala 34:12]
  wire [31:0] _GEN_657; // @[FFT.scala 34:12]
  wire [31:0] _GEN_658; // @[FFT.scala 34:12]
  wire [31:0] _GEN_659; // @[FFT.scala 34:12]
  wire [31:0] _GEN_660; // @[FFT.scala 34:12]
  wire [31:0] _GEN_661; // @[FFT.scala 34:12]
  wire [31:0] _GEN_662; // @[FFT.scala 34:12]
  wire [31:0] _GEN_663; // @[FFT.scala 34:12]
  wire [31:0] _GEN_664; // @[FFT.scala 34:12]
  wire [31:0] _GEN_665; // @[FFT.scala 34:12]
  wire [31:0] _GEN_666; // @[FFT.scala 34:12]
  wire [31:0] _GEN_667; // @[FFT.scala 34:12]
  wire [31:0] _GEN_668; // @[FFT.scala 34:12]
  wire [31:0] _GEN_669; // @[FFT.scala 34:12]
  wire [31:0] _GEN_670; // @[FFT.scala 34:12]
  wire [31:0] _GEN_671; // @[FFT.scala 34:12]
  wire [31:0] _GEN_672; // @[FFT.scala 34:12]
  wire [31:0] _GEN_673; // @[FFT.scala 34:12]
  wire [31:0] _GEN_674; // @[FFT.scala 34:12]
  wire [31:0] _GEN_675; // @[FFT.scala 34:12]
  wire [31:0] _GEN_676; // @[FFT.scala 34:12]
  wire [31:0] _GEN_677; // @[FFT.scala 34:12]
  wire [31:0] _GEN_678; // @[FFT.scala 34:12]
  wire [31:0] _GEN_679; // @[FFT.scala 34:12]
  wire [31:0] _GEN_680; // @[FFT.scala 34:12]
  wire [31:0] _GEN_681; // @[FFT.scala 34:12]
  wire [31:0] _GEN_682; // @[FFT.scala 34:12]
  wire [31:0] _GEN_683; // @[FFT.scala 34:12]
  wire [31:0] _GEN_684; // @[FFT.scala 34:12]
  wire [31:0] _GEN_685; // @[FFT.scala 34:12]
  wire [31:0] _GEN_686; // @[FFT.scala 34:12]
  wire [31:0] _GEN_687; // @[FFT.scala 34:12]
  wire [31:0] _GEN_688; // @[FFT.scala 34:12]
  wire [31:0] _GEN_689; // @[FFT.scala 34:12]
  wire [31:0] _GEN_690; // @[FFT.scala 34:12]
  wire [31:0] _GEN_691; // @[FFT.scala 34:12]
  wire [31:0] _GEN_692; // @[FFT.scala 34:12]
  wire [31:0] _GEN_693; // @[FFT.scala 34:12]
  wire [31:0] _GEN_694; // @[FFT.scala 34:12]
  wire [31:0] _GEN_695; // @[FFT.scala 34:12]
  wire [31:0] _GEN_696; // @[FFT.scala 34:12]
  wire [31:0] _GEN_697; // @[FFT.scala 34:12]
  wire [31:0] _GEN_698; // @[FFT.scala 34:12]
  wire [31:0] _GEN_699; // @[FFT.scala 34:12]
  wire [31:0] _GEN_700; // @[FFT.scala 34:12]
  wire [31:0] _GEN_701; // @[FFT.scala 34:12]
  wire [31:0] _GEN_702; // @[FFT.scala 34:12]
  wire [31:0] _GEN_703; // @[FFT.scala 34:12]
  wire [31:0] _GEN_706; // @[FFT.scala 35:12]
  wire [31:0] _GEN_707; // @[FFT.scala 35:12]
  wire [31:0] _GEN_708; // @[FFT.scala 35:12]
  wire [31:0] _GEN_709; // @[FFT.scala 35:12]
  wire [31:0] _GEN_710; // @[FFT.scala 35:12]
  wire [31:0] _GEN_711; // @[FFT.scala 35:12]
  wire [31:0] _GEN_712; // @[FFT.scala 35:12]
  wire [31:0] _GEN_713; // @[FFT.scala 35:12]
  wire [31:0] _GEN_714; // @[FFT.scala 35:12]
  wire [31:0] _GEN_715; // @[FFT.scala 35:12]
  wire [31:0] _GEN_716; // @[FFT.scala 35:12]
  wire [31:0] _GEN_717; // @[FFT.scala 35:12]
  wire [31:0] _GEN_718; // @[FFT.scala 35:12]
  wire [31:0] _GEN_719; // @[FFT.scala 35:12]
  wire [31:0] _GEN_720; // @[FFT.scala 35:12]
  wire [31:0] _GEN_721; // @[FFT.scala 35:12]
  wire [31:0] _GEN_722; // @[FFT.scala 35:12]
  wire [31:0] _GEN_723; // @[FFT.scala 35:12]
  wire [31:0] _GEN_724; // @[FFT.scala 35:12]
  wire [31:0] _GEN_725; // @[FFT.scala 35:12]
  wire [31:0] _GEN_726; // @[FFT.scala 35:12]
  wire [31:0] _GEN_727; // @[FFT.scala 35:12]
  wire [31:0] _GEN_728; // @[FFT.scala 35:12]
  wire [31:0] _GEN_729; // @[FFT.scala 35:12]
  wire [31:0] _GEN_730; // @[FFT.scala 35:12]
  wire [31:0] _GEN_731; // @[FFT.scala 35:12]
  wire [31:0] _GEN_732; // @[FFT.scala 35:12]
  wire [31:0] _GEN_733; // @[FFT.scala 35:12]
  wire [31:0] _GEN_734; // @[FFT.scala 35:12]
  wire [31:0] _GEN_735; // @[FFT.scala 35:12]
  wire [31:0] _GEN_736; // @[FFT.scala 35:12]
  wire [31:0] _GEN_737; // @[FFT.scala 35:12]
  wire [31:0] _GEN_738; // @[FFT.scala 35:12]
  wire [31:0] _GEN_739; // @[FFT.scala 35:12]
  wire [31:0] _GEN_740; // @[FFT.scala 35:12]
  wire [31:0] _GEN_741; // @[FFT.scala 35:12]
  wire [31:0] _GEN_742; // @[FFT.scala 35:12]
  wire [31:0] _GEN_743; // @[FFT.scala 35:12]
  wire [31:0] _GEN_744; // @[FFT.scala 35:12]
  wire [31:0] _GEN_745; // @[FFT.scala 35:12]
  wire [31:0] _GEN_746; // @[FFT.scala 35:12]
  wire [31:0] _GEN_747; // @[FFT.scala 35:12]
  wire [31:0] _GEN_748; // @[FFT.scala 35:12]
  wire [31:0] _GEN_749; // @[FFT.scala 35:12]
  wire [31:0] _GEN_750; // @[FFT.scala 35:12]
  wire [31:0] _GEN_751; // @[FFT.scala 35:12]
  wire [31:0] _GEN_752; // @[FFT.scala 35:12]
  wire [31:0] _GEN_753; // @[FFT.scala 35:12]
  wire [31:0] _GEN_754; // @[FFT.scala 35:12]
  wire [31:0] _GEN_755; // @[FFT.scala 35:12]
  wire [31:0] _GEN_756; // @[FFT.scala 35:12]
  wire [31:0] _GEN_757; // @[FFT.scala 35:12]
  wire [31:0] _GEN_758; // @[FFT.scala 35:12]
  wire [31:0] _GEN_759; // @[FFT.scala 35:12]
  wire [31:0] _GEN_760; // @[FFT.scala 35:12]
  wire [31:0] _GEN_761; // @[FFT.scala 35:12]
  wire [31:0] _GEN_762; // @[FFT.scala 35:12]
  wire [31:0] _GEN_763; // @[FFT.scala 35:12]
  wire [31:0] _GEN_764; // @[FFT.scala 35:12]
  wire [31:0] _GEN_765; // @[FFT.scala 35:12]
  wire [31:0] _GEN_766; // @[FFT.scala 35:12]
  wire [31:0] _GEN_767; // @[FFT.scala 35:12]
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_521;
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_522;
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_523;
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_524;
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_525;
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_526;
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_527;
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_528;
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_529;
  reg [31:0] _T_402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_530;
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_531;
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_532;
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_533;
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_534;
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_535;
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_536;
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_537;
  reg [31:0] _T_406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_538;
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_539;
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_540;
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_541;
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [31:0] _T_409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  reg [31:0] _T_409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_552;
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_553;
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_554;
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_557;
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_558;
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_559;
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_560;
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_561;
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_562;
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_563;
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_564;
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_565;
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_566;
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_567;
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_568;
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_569;
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_570;
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_571;
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_572;
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_573;
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_574;
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_575;
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_576;
  wire [31:0] _GEN_962; // @[FFT.scala 34:12]
  wire [31:0] _GEN_963; // @[FFT.scala 34:12]
  wire [31:0] _GEN_964; // @[FFT.scala 34:12]
  wire [31:0] _GEN_965; // @[FFT.scala 34:12]
  wire [31:0] _GEN_966; // @[FFT.scala 34:12]
  wire [31:0] _GEN_967; // @[FFT.scala 34:12]
  wire [31:0] _GEN_968; // @[FFT.scala 34:12]
  wire [31:0] _GEN_969; // @[FFT.scala 34:12]
  wire [31:0] _GEN_970; // @[FFT.scala 34:12]
  wire [31:0] _GEN_971; // @[FFT.scala 34:12]
  wire [31:0] _GEN_972; // @[FFT.scala 34:12]
  wire [31:0] _GEN_973; // @[FFT.scala 34:12]
  wire [31:0] _GEN_974; // @[FFT.scala 34:12]
  wire [31:0] _GEN_975; // @[FFT.scala 34:12]
  wire [31:0] _GEN_976; // @[FFT.scala 34:12]
  wire [31:0] _GEN_977; // @[FFT.scala 34:12]
  wire [31:0] _GEN_978; // @[FFT.scala 34:12]
  wire [31:0] _GEN_979; // @[FFT.scala 34:12]
  wire [31:0] _GEN_980; // @[FFT.scala 34:12]
  wire [31:0] _GEN_981; // @[FFT.scala 34:12]
  wire [31:0] _GEN_982; // @[FFT.scala 34:12]
  wire [31:0] _GEN_983; // @[FFT.scala 34:12]
  wire [31:0] _GEN_984; // @[FFT.scala 34:12]
  wire [31:0] _GEN_985; // @[FFT.scala 34:12]
  wire [31:0] _GEN_986; // @[FFT.scala 34:12]
  wire [31:0] _GEN_987; // @[FFT.scala 34:12]
  wire [31:0] _GEN_988; // @[FFT.scala 34:12]
  wire [31:0] _GEN_989; // @[FFT.scala 34:12]
  wire [31:0] _GEN_990; // @[FFT.scala 34:12]
  wire [31:0] _GEN_991; // @[FFT.scala 34:12]
  wire [31:0] _GEN_994; // @[FFT.scala 35:12]
  wire [31:0] _GEN_995; // @[FFT.scala 35:12]
  wire [31:0] _GEN_996; // @[FFT.scala 35:12]
  wire [31:0] _GEN_997; // @[FFT.scala 35:12]
  wire [31:0] _GEN_998; // @[FFT.scala 35:12]
  wire [31:0] _GEN_999; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1000; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1001; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1002; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1003; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1004; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1005; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1006; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1007; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1008; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1009; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1010; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1011; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1012; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1013; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1014; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1015; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1016; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1017; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1018; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1019; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1020; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1021; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1022; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1023; // @[FFT.scala 35:12]
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_577;
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_578;
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_579;
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_580;
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_581;
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_582;
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_583;
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_584;
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_585;
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_586;
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_587;
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_588;
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_589;
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_590;
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_591;
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_592;
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_593;
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_594;
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_595;
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_596;
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_597;
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_598;
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_599;
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_600;
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_601;
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_602;
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_603;
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_604;
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_605;
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_606;
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_607;
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_608;
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_609;
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_610;
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_611;
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_612;
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_613;
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_614;
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_615;
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_616;
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_617;
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_618;
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_619;
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_620;
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_621;
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_622;
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_623;
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_624;
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_625;
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_626;
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_627;
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_628;
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_629;
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_630;
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_631;
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_632;
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_633;
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_634;
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_635;
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_636;
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_637;
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_638;
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_639;
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_640;
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_641;
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_642;
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_643;
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_644;
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_645;
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_646;
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_647;
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_648;
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_649;
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_650;
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_651;
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_652;
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_653;
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_654;
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_655;
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_656;
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_657;
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_658;
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_659;
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_660;
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_661;
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_662;
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_663;
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_664;
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_665;
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_666;
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_667;
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_668;
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_669;
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_670;
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_671;
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_672;
  wire [31:0] _GEN_1122; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1123; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1124; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1125; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1126; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1127; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1128; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1129; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1130; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1131; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1132; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1133; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1134; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1135; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1138; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1139; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1140; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1141; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1142; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1143; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1144; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1145; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1146; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1147; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1148; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1149; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1150; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1151; // @[FFT.scala 35:12]
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_673;
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_674;
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_675;
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_676;
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_677;
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_678;
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_679;
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_680;
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_681;
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_682;
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_683;
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_684;
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_685;
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_686;
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_687;
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_688;
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_689;
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_690;
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_691;
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_692;
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_693;
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_694;
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_695;
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_696;
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_697;
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_698;
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_699;
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_700;
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_701;
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_702;
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_703;
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_704;
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_705;
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_706;
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_707;
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_708;
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_709;
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_710;
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_711;
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_712;
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_713;
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_714;
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_715;
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_716;
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_717;
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_718;
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_719;
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_720;
  wire [31:0] _GEN_1202; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1203; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1204; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1205; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1206; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1207; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1210; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1211; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1212; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1213; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1214; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1215; // @[FFT.scala 35:12]
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_721;
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_722;
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_723;
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_724;
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_725;
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_726;
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_727;
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_728;
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_729;
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_730;
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_731;
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_732;
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_733;
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_734;
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_735;
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_736;
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_737;
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_738;
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_739;
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_740;
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_741;
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_742;
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_743;
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_744;
  wire [31:0] _GEN_1242; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1243; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1246; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1247; // @[FFT.scala 35:12]
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_745;
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_746;
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_747;
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_748;
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_749;
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_750;
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_751;
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_752;
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_753;
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_754;
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_755;
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_756;
  reg [31:0] _T_540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_757;
  reg [31:0] _T_540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_758;
  reg [31:0] _T_541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_759;
  reg [31:0] _T_541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_760;
  reg [31:0] _T_543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_761;
  reg [31:0] _T_543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_762;
  reg [31:0] out1D1_re; // @[FFT.scala 58:23]
  reg [31:0] _RAND_763;
  reg [31:0] out1D1_im; // @[FFT.scala 58:23]
  reg [31:0] _RAND_764;
  reg [31:0] _T_544_re; // @[FFT.scala 62:22]
  reg [31:0] _RAND_765;
  reg [31:0] _T_544_im; // @[FFT.scala 62:22]
  reg [31:0] _RAND_766;
  reg [31:0] _T_545_re; // @[FFT.scala 63:22]
  reg [31:0] _RAND_767;
  reg [31:0] _T_545_im; // @[FFT.scala 63:22]
  reg [31:0] _RAND_768;
  reg  _T_546; // @[Reg.scala 15:16]
  reg [31:0] _RAND_769;
  reg  _T_547; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  reg  _T_548; // @[Reg.scala 15:16]
  reg [31:0] _RAND_771;
  reg  _T_549; // @[Reg.scala 15:16]
  reg [31:0] _RAND_772;
  reg  _T_550; // @[Reg.scala 15:16]
  reg [31:0] _RAND_773;
  reg  _T_551; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  reg  _T_552; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  reg  _T_553; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  reg  _T_554; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg  _T_555; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  reg  _T_556; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg  _T_557; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  reg  _T_558; // @[Reg.scala 15:16]
  reg [31:0] _RAND_781;
  reg  _T_559; // @[Reg.scala 15:16]
  reg [31:0] _RAND_782;
  reg  _T_560; // @[Reg.scala 15:16]
  reg [31:0] _RAND_783;
  reg  _T_561; // @[Reg.scala 15:16]
  reg [31:0] _RAND_784;
  reg  _T_562; // @[Reg.scala 15:16]
  reg [31:0] _RAND_785;
  reg  _T_563; // @[Reg.scala 15:16]
  reg [31:0] _RAND_786;
  reg  _T_564; // @[Reg.scala 15:16]
  reg [31:0] _RAND_787;
  reg  _T_565; // @[Reg.scala 15:16]
  reg [31:0] _RAND_788;
  reg  _T_566; // @[Reg.scala 15:16]
  reg [31:0] _RAND_789;
  reg  _T_567; // @[Reg.scala 15:16]
  reg [31:0] _RAND_790;
  reg  _T_568; // @[Reg.scala 15:16]
  reg [31:0] _RAND_791;
  reg  _T_569; // @[Reg.scala 15:16]
  reg [31:0] _RAND_792;
  reg  _T_570; // @[Reg.scala 15:16]
  reg [31:0] _RAND_793;
  reg  _T_571; // @[Reg.scala 15:16]
  reg [31:0] _RAND_794;
  reg  _T_572; // @[Reg.scala 15:16]
  reg [31:0] _RAND_795;
  reg  _T_573; // @[Reg.scala 15:16]
  reg [31:0] _RAND_796;
  reg  _T_574; // @[Reg.scala 15:16]
  reg [31:0] _RAND_797;
  reg  _T_575; // @[Reg.scala 15:16]
  reg [31:0] _RAND_798;
  reg  _T_576; // @[Reg.scala 15:16]
  reg [31:0] _RAND_799;
  reg  _T_577; // @[Reg.scala 15:16]
  reg [31:0] _RAND_800;
  reg  _T_578; // @[Reg.scala 15:16]
  reg [31:0] _RAND_801;
  reg  _T_579; // @[Reg.scala 15:16]
  reg [31:0] _RAND_802;
  reg  _T_580; // @[Reg.scala 15:16]
  reg [31:0] _RAND_803;
  reg  _T_581; // @[Reg.scala 15:16]
  reg [31:0] _RAND_804;
  reg  _T_582; // @[Reg.scala 15:16]
  reg [31:0] _RAND_805;
  reg  _T_583; // @[Reg.scala 15:16]
  reg [31:0] _RAND_806;
  reg  _T_584; // @[Reg.scala 15:16]
  reg [31:0] _RAND_807;
  reg  _T_585; // @[Reg.scala 15:16]
  reg [31:0] _RAND_808;
  reg  _T_586; // @[Reg.scala 15:16]
  reg [31:0] _RAND_809;
  reg  _T_587; // @[Reg.scala 15:16]
  reg [31:0] _RAND_810;
  reg  _T_588; // @[Reg.scala 15:16]
  reg [31:0] _RAND_811;
  reg  _T_589; // @[Reg.scala 15:16]
  reg [31:0] _RAND_812;
  reg  _T_590; // @[Reg.scala 15:16]
  reg [31:0] _RAND_813;
  reg  _T_591; // @[Reg.scala 15:16]
  reg [31:0] _RAND_814;
  reg  _T_592; // @[Reg.scala 15:16]
  reg [31:0] _RAND_815;
  reg  _T_593; // @[Reg.scala 15:16]
  reg [31:0] _RAND_816;
  reg  _T_594; // @[Reg.scala 15:16]
  reg [31:0] _RAND_817;
  reg  _T_595; // @[Reg.scala 15:16]
  reg [31:0] _RAND_818;
  reg  _T_596; // @[Reg.scala 15:16]
  reg [31:0] _RAND_819;
  reg  _T_597; // @[Reg.scala 15:16]
  reg [31:0] _RAND_820;
  reg  _T_598; // @[Reg.scala 15:16]
  reg [31:0] _RAND_821;
  reg  _T_599; // @[Reg.scala 15:16]
  reg [31:0] _RAND_822;
  reg  _T_600; // @[Reg.scala 15:16]
  reg [31:0] _RAND_823;
  reg  _T_601; // @[Reg.scala 15:16]
  reg [31:0] _RAND_824;
  reg  _T_602; // @[Reg.scala 15:16]
  reg [31:0] _RAND_825;
  reg  _T_603; // @[Reg.scala 15:16]
  reg [31:0] _RAND_826;
  reg  _T_604; // @[Reg.scala 15:16]
  reg [31:0] _RAND_827;
  reg  _T_605; // @[Reg.scala 15:16]
  reg [31:0] _RAND_828;
  reg  _T_606; // @[Reg.scala 15:16]
  reg [31:0] _RAND_829;
  reg  _T_607; // @[Reg.scala 15:16]
  reg [31:0] _RAND_830;
  reg  _T_608; // @[Reg.scala 15:16]
  reg [31:0] _RAND_831;
  reg  _T_609; // @[Reg.scala 15:16]
  reg [31:0] _RAND_832;
  reg  _T_610; // @[Reg.scala 15:16]
  reg [31:0] _RAND_833;
  reg  _T_611; // @[Reg.scala 15:16]
  reg [31:0] _RAND_834;
  reg  _T_612; // @[Reg.scala 15:16]
  reg [31:0] _RAND_835;
  reg  _T_613; // @[Reg.scala 15:16]
  reg [31:0] _RAND_836;
  reg  _T_614; // @[Reg.scala 15:16]
  reg [31:0] _RAND_837;
  reg  _T_615; // @[Reg.scala 15:16]
  reg [31:0] _RAND_838;
  reg  _T_616; // @[Reg.scala 15:16]
  reg [31:0] _RAND_839;
  reg  _T_617; // @[Reg.scala 15:16]
  reg [31:0] _RAND_840;
  reg  _T_618; // @[Reg.scala 15:16]
  reg [31:0] _RAND_841;
  reg  _T_619; // @[Reg.scala 15:16]
  reg [31:0] _RAND_842;
  reg  _T_620; // @[Reg.scala 15:16]
  reg [31:0] _RAND_843;
  reg  _T_621; // @[Reg.scala 15:16]
  reg [31:0] _RAND_844;
  reg  _T_622; // @[Reg.scala 15:16]
  reg [31:0] _RAND_845;
  reg  _T_623; // @[Reg.scala 15:16]
  reg [31:0] _RAND_846;
  reg  _T_624; // @[Reg.scala 15:16]
  reg [31:0] _RAND_847;
  reg  _T_625; // @[Reg.scala 15:16]
  reg [31:0] _RAND_848;
  reg  _T_626; // @[Reg.scala 15:16]
  reg [31:0] _RAND_849;
  reg  _T_627; // @[Reg.scala 15:16]
  reg [31:0] _RAND_850;
  reg  _T_628; // @[Reg.scala 15:16]
  reg [31:0] _RAND_851;
  reg  _T_629; // @[Reg.scala 15:16]
  reg [31:0] _RAND_852;
  reg  _T_630; // @[Reg.scala 15:16]
  reg [31:0] _RAND_853;
  reg  _T_631; // @[Reg.scala 15:16]
  reg [31:0] _RAND_854;
  reg  _T_632; // @[Reg.scala 15:16]
  reg [31:0] _RAND_855;
  reg  _T_633; // @[Reg.scala 15:16]
  reg [31:0] _RAND_856;
  reg  _T_634; // @[Reg.scala 15:16]
  reg [31:0] _RAND_857;
  reg  _T_635; // @[Reg.scala 15:16]
  reg [31:0] _RAND_858;
  reg  _T_636; // @[Reg.scala 15:16]
  reg [31:0] _RAND_859;
  reg  _T_637; // @[Reg.scala 15:16]
  reg [31:0] _RAND_860;
  reg  _T_638; // @[Reg.scala 15:16]
  reg [31:0] _RAND_861;
  reg  _T_639; // @[Reg.scala 15:16]
  reg [31:0] _RAND_862;
  reg  _T_640; // @[Reg.scala 15:16]
  reg [31:0] _RAND_863;
  reg  _T_641; // @[Reg.scala 15:16]
  reg [31:0] _RAND_864;
  reg  _T_642; // @[Reg.scala 15:16]
  reg [31:0] _RAND_865;
  reg  _T_643; // @[Reg.scala 15:16]
  reg [31:0] _RAND_866;
  reg  _T_644; // @[Reg.scala 15:16]
  reg [31:0] _RAND_867;
  reg  _T_645; // @[Reg.scala 15:16]
  reg [31:0] _RAND_868;
  reg  _T_646; // @[Reg.scala 15:16]
  reg [31:0] _RAND_869;
  reg  _T_647; // @[Reg.scala 15:16]
  reg [31:0] _RAND_870;
  reg  _T_648; // @[Reg.scala 15:16]
  reg [31:0] _RAND_871;
  reg  _T_649; // @[Reg.scala 15:16]
  reg [31:0] _RAND_872;
  reg  _T_650; // @[Reg.scala 15:16]
  reg [31:0] _RAND_873;
  reg  _T_651; // @[Reg.scala 15:16]
  reg [31:0] _RAND_874;
  reg  _T_652; // @[Reg.scala 15:16]
  reg [31:0] _RAND_875;
  reg  _T_653; // @[Reg.scala 15:16]
  reg [31:0] _RAND_876;
  reg  _T_654; // @[Reg.scala 15:16]
  reg [31:0] _RAND_877;
  reg  _T_655; // @[Reg.scala 15:16]
  reg [31:0] _RAND_878;
  reg  _T_656; // @[Reg.scala 15:16]
  reg [31:0] _RAND_879;
  reg  _T_657; // @[Reg.scala 15:16]
  reg [31:0] _RAND_880;
  reg  _T_658; // @[Reg.scala 15:16]
  reg [31:0] _RAND_881;
  reg  _T_659; // @[Reg.scala 15:16]
  reg [31:0] _RAND_882;
  reg  _T_660; // @[Reg.scala 15:16]
  reg [31:0] _RAND_883;
  reg  _T_661; // @[Reg.scala 15:16]
  reg [31:0] _RAND_884;
  reg  _T_662; // @[Reg.scala 15:16]
  reg [31:0] _RAND_885;
  reg  _T_663; // @[Reg.scala 15:16]
  reg [31:0] _RAND_886;
  reg  _T_664; // @[Reg.scala 15:16]
  reg [31:0] _RAND_887;
  reg  _T_665; // @[Reg.scala 15:16]
  reg [31:0] _RAND_888;
  reg  _T_666; // @[Reg.scala 15:16]
  reg [31:0] _RAND_889;
  reg  _T_667; // @[Reg.scala 15:16]
  reg [31:0] _RAND_890;
  reg  _T_668; // @[Reg.scala 15:16]
  reg [31:0] _RAND_891;
  reg  _T_669; // @[Reg.scala 15:16]
  reg [31:0] _RAND_892;
  reg  _T_670; // @[Reg.scala 15:16]
  reg [31:0] _RAND_893;
  reg  _T_671; // @[Reg.scala 15:16]
  reg [31:0] _RAND_894;
  reg  _T_672; // @[Reg.scala 15:16]
  reg [31:0] _RAND_895;
  reg  _T_673; // @[Reg.scala 15:16]
  reg [31:0] _RAND_896;
  reg  _T_674; // @[Reg.scala 15:16]
  reg [31:0] _RAND_897;
  reg  _T_675; // @[Reg.scala 15:16]
  reg [31:0] _RAND_898;
  reg  _T_676; // @[Reg.scala 15:16]
  reg [31:0] _RAND_899;
  reg  _T_677; // @[Reg.scala 15:16]
  reg [31:0] _RAND_900;
  reg  _T_678; // @[Reg.scala 15:16]
  reg [31:0] _RAND_901;
  reg  _T_679; // @[Reg.scala 15:16]
  reg [31:0] _RAND_902;
  reg  _T_680; // @[Reg.scala 15:16]
  reg [31:0] _RAND_903;
  reg  _T_681; // @[Reg.scala 15:16]
  reg [31:0] _RAND_904;
  reg  _T_682; // @[Reg.scala 15:16]
  reg [31:0] _RAND_905;
  reg  _T_683; // @[Reg.scala 15:16]
  reg [31:0] _RAND_906;
  reg  _T_684; // @[Reg.scala 15:16]
  reg [31:0] _RAND_907;
  reg  _T_685; // @[Reg.scala 15:16]
  reg [31:0] _RAND_908;
  reg  _T_686; // @[Reg.scala 15:16]
  reg [31:0] _RAND_909;
  reg  _T_687; // @[Reg.scala 15:16]
  reg [31:0] _RAND_910;
  reg  _T_688; // @[Reg.scala 15:16]
  reg [31:0] _RAND_911;
  reg  _T_689; // @[Reg.scala 15:16]
  reg [31:0] _RAND_912;
  reg  _T_690; // @[Reg.scala 15:16]
  reg [31:0] _RAND_913;
  reg  _T_691; // @[Reg.scala 15:16]
  reg [31:0] _RAND_914;
  reg  _T_692; // @[Reg.scala 15:16]
  reg [31:0] _RAND_915;
  reg  _T_693; // @[Reg.scala 15:16]
  reg [31:0] _RAND_916;
  reg  _T_694; // @[Reg.scala 15:16]
  reg [31:0] _RAND_917;
  reg  _T_695; // @[Reg.scala 15:16]
  reg [31:0] _RAND_918;
  reg  _T_696; // @[Reg.scala 15:16]
  reg [31:0] _RAND_919;
  reg  _T_697; // @[Reg.scala 15:16]
  reg [31:0] _RAND_920;
  reg  _T_698; // @[Reg.scala 15:16]
  reg [31:0] _RAND_921;
  reg  _T_699; // @[Reg.scala 15:16]
  reg [31:0] _RAND_922;
  reg  _T_700; // @[Reg.scala 15:16]
  reg [31:0] _RAND_923;
  reg  _T_701; // @[Reg.scala 15:16]
  reg [31:0] _RAND_924;
  reg  _T_702; // @[Reg.scala 15:16]
  reg [31:0] _RAND_925;
  reg  _T_703; // @[Reg.scala 15:16]
  reg [31:0] _RAND_926;
  reg  _T_704; // @[Reg.scala 15:16]
  reg [31:0] _RAND_927;
  reg  _T_705; // @[Reg.scala 15:16]
  reg [31:0] _RAND_928;
  reg  _T_706; // @[Reg.scala 15:16]
  reg [31:0] _RAND_929;
  reg  _T_707; // @[Reg.scala 15:16]
  reg [31:0] _RAND_930;
  reg  _T_708; // @[Reg.scala 15:16]
  reg [31:0] _RAND_931;
  reg  _T_709; // @[Reg.scala 15:16]
  reg [31:0] _RAND_932;
  reg  _T_710; // @[Reg.scala 15:16]
  reg [31:0] _RAND_933;
  reg  _T_711; // @[Reg.scala 15:16]
  reg [31:0] _RAND_934;
  reg  _T_712; // @[Reg.scala 15:16]
  reg [31:0] _RAND_935;
  reg  _T_713; // @[Reg.scala 15:16]
  reg [31:0] _RAND_936;
  reg  _T_714; // @[Reg.scala 15:16]
  reg [31:0] _RAND_937;
  reg  _T_715; // @[Reg.scala 15:16]
  reg [31:0] _RAND_938;
  reg  _T_716; // @[Reg.scala 15:16]
  reg [31:0] _RAND_939;
  reg  _T_717; // @[Reg.scala 15:16]
  reg [31:0] _RAND_940;
  reg  _T_718; // @[Reg.scala 15:16]
  reg [31:0] _RAND_941;
  reg  _T_719; // @[Reg.scala 15:16]
  reg [31:0] _RAND_942;
  reg  _T_720; // @[Reg.scala 15:16]
  reg [31:0] _RAND_943;
  reg  _T_721; // @[Reg.scala 15:16]
  reg [31:0] _RAND_944;
  reg  _T_722; // @[Reg.scala 15:16]
  reg [31:0] _RAND_945;
  reg  _T_723; // @[Reg.scala 15:16]
  reg [31:0] _RAND_946;
  reg  _T_724; // @[Reg.scala 15:16]
  reg [31:0] _RAND_947;
  reg  _T_725; // @[Reg.scala 15:16]
  reg [31:0] _RAND_948;
  reg  _T_726; // @[Reg.scala 15:16]
  reg [31:0] _RAND_949;
  reg  _T_727; // @[Reg.scala 15:16]
  reg [31:0] _RAND_950;
  reg  _T_728; // @[Reg.scala 15:16]
  reg [31:0] _RAND_951;
  reg  _T_729; // @[Reg.scala 15:16]
  reg [31:0] _RAND_952;
  reg  _T_730; // @[Reg.scala 15:16]
  reg [31:0] _RAND_953;
  reg  _T_731; // @[Reg.scala 15:16]
  reg [31:0] _RAND_954;
  reg  _T_732; // @[Reg.scala 15:16]
  reg [31:0] _RAND_955;
  reg  _T_733; // @[Reg.scala 15:16]
  reg [31:0] _RAND_956;
  reg  _T_734; // @[Reg.scala 15:16]
  reg [31:0] _RAND_957;
  reg  _T_735; // @[Reg.scala 15:16]
  reg [31:0] _RAND_958;
  reg  _T_736; // @[Reg.scala 15:16]
  reg [31:0] _RAND_959;
  reg  _T_737; // @[Reg.scala 15:16]
  reg [31:0] _RAND_960;
  reg  _T_738; // @[Reg.scala 15:16]
  reg [31:0] _RAND_961;
  reg  _T_739; // @[Reg.scala 15:16]
  reg [31:0] _RAND_962;
  reg  _T_740; // @[Reg.scala 15:16]
  reg [31:0] _RAND_963;
  reg  _T_741; // @[Reg.scala 15:16]
  reg [31:0] _RAND_964;
  reg  _T_742; // @[Reg.scala 15:16]
  reg [31:0] _RAND_965;
  reg  _T_743; // @[Reg.scala 15:16]
  reg [31:0] _RAND_966;
  reg  _T_744; // @[Reg.scala 15:16]
  reg [31:0] _RAND_967;
  reg  _T_745; // @[Reg.scala 15:16]
  reg [31:0] _RAND_968;
  reg  _T_746; // @[Reg.scala 15:16]
  reg [31:0] _RAND_969;
  reg  _T_747; // @[Reg.scala 15:16]
  reg [31:0] _RAND_970;
  reg  _T_748; // @[Reg.scala 15:16]
  reg [31:0] _RAND_971;
  reg  _T_749; // @[Reg.scala 15:16]
  reg [31:0] _RAND_972;
  reg  _T_750; // @[Reg.scala 15:16]
  reg [31:0] _RAND_973;
  reg  _T_751; // @[Reg.scala 15:16]
  reg [31:0] _RAND_974;
  reg  _T_752; // @[Reg.scala 15:16]
  reg [31:0] _RAND_975;
  reg  _T_753; // @[Reg.scala 15:16]
  reg [31:0] _RAND_976;
  reg  _T_754; // @[Reg.scala 15:16]
  reg [31:0] _RAND_977;
  reg  _T_755; // @[Reg.scala 15:16]
  reg [31:0] _RAND_978;
  reg  _T_756; // @[Reg.scala 15:16]
  reg [31:0] _RAND_979;
  reg  _T_757; // @[Reg.scala 15:16]
  reg [31:0] _RAND_980;
  reg  _T_758; // @[Reg.scala 15:16]
  reg [31:0] _RAND_981;
  reg  _T_759; // @[Reg.scala 15:16]
  reg [31:0] _RAND_982;
  reg  _T_760; // @[Reg.scala 15:16]
  reg [31:0] _RAND_983;
  reg  _T_761; // @[Reg.scala 15:16]
  reg [31:0] _RAND_984;
  reg  _T_762; // @[Reg.scala 15:16]
  reg [31:0] _RAND_985;
  reg  _T_763; // @[Reg.scala 15:16]
  reg [31:0] _RAND_986;
  reg  _T_764; // @[Reg.scala 15:16]
  reg [31:0] _RAND_987;
  reg  _T_765; // @[Reg.scala 15:16]
  reg [31:0] _RAND_988;
  reg  _T_766; // @[Reg.scala 15:16]
  reg [31:0] _RAND_989;
  reg  _T_767; // @[Reg.scala 15:16]
  reg [31:0] _RAND_990;
  reg  _T_768; // @[Reg.scala 15:16]
  reg [31:0] _RAND_991;
  reg  _T_769; // @[Reg.scala 15:16]
  reg [31:0] _RAND_992;
  reg  _T_770; // @[Reg.scala 15:16]
  reg [31:0] _RAND_993;
  reg  _T_771; // @[Reg.scala 15:16]
  reg [31:0] _RAND_994;
  reg  _T_772; // @[Reg.scala 15:16]
  reg [31:0] _RAND_995;
  reg  _T_773; // @[Reg.scala 15:16]
  reg [31:0] _RAND_996;
  reg  _T_774; // @[Reg.scala 15:16]
  reg [31:0] _RAND_997;
  reg  _T_775; // @[Reg.scala 15:16]
  reg [31:0] _RAND_998;
  reg  _T_776; // @[Reg.scala 15:16]
  reg [31:0] _RAND_999;
  reg  _T_777; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1000;
  reg  _T_778; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1001;
  reg  _T_779; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1002;
  reg  _T_780; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1003;
  reg  _T_781; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1004;
  reg  _T_782; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1005;
  reg  _T_783; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1006;
  reg  _T_784; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1007;
  reg  _T_785; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1008;
  reg  _T_786; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1009;
  reg  _T_787; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1010;
  reg  _T_788; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1011;
  reg  _T_789; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1012;
  reg  _T_790; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1013;
  reg  _T_791; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1014;
  reg  _T_792; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1015;
  reg  _T_793; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1016;
  reg  _T_794; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1017;
  reg  _T_795; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1018;
  reg  _T_796; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1019;
  reg  _T_797; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1020;
  reg  _T_798; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1021;
  reg  _T_799; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1022;
  reg  _T_800; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1023;
  reg  _T_801; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1024;
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign _T_1 = cnt + 8'h1; // @[FFT.scala 42:16]
  assign _GEN_2 = 7'h1 == cnt[6:0] ? $signed(32'shffec) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_3 = 7'h2 == cnt[6:0] ? $signed(32'shffb1) : $signed(_GEN_2); // @[FFT.scala 34:12]
  assign _GEN_4 = 7'h3 == cnt[6:0] ? $signed(32'shff4e) : $signed(_GEN_3); // @[FFT.scala 34:12]
  assign _GEN_5 = 7'h4 == cnt[6:0] ? $signed(32'shfec4) : $signed(_GEN_4); // @[FFT.scala 34:12]
  assign _GEN_6 = 7'h5 == cnt[6:0] ? $signed(32'shfe13) : $signed(_GEN_5); // @[FFT.scala 34:12]
  assign _GEN_7 = 7'h6 == cnt[6:0] ? $signed(32'shfd3b) : $signed(_GEN_6); // @[FFT.scala 34:12]
  assign _GEN_8 = 7'h7 == cnt[6:0] ? $signed(32'shfc3b) : $signed(_GEN_7); // @[FFT.scala 34:12]
  assign _GEN_9 = 7'h8 == cnt[6:0] ? $signed(32'shfb15) : $signed(_GEN_8); // @[FFT.scala 34:12]
  assign _GEN_10 = 7'h9 == cnt[6:0] ? $signed(32'shf9c8) : $signed(_GEN_9); // @[FFT.scala 34:12]
  assign _GEN_11 = 7'ha == cnt[6:0] ? $signed(32'shf854) : $signed(_GEN_10); // @[FFT.scala 34:12]
  assign _GEN_12 = 7'hb == cnt[6:0] ? $signed(32'shf6ba) : $signed(_GEN_11); // @[FFT.scala 34:12]
  assign _GEN_13 = 7'hc == cnt[6:0] ? $signed(32'shf4fa) : $signed(_GEN_12); // @[FFT.scala 34:12]
  assign _GEN_14 = 7'hd == cnt[6:0] ? $signed(32'shf314) : $signed(_GEN_13); // @[FFT.scala 34:12]
  assign _GEN_15 = 7'he == cnt[6:0] ? $signed(32'shf109) : $signed(_GEN_14); // @[FFT.scala 34:12]
  assign _GEN_16 = 7'hf == cnt[6:0] ? $signed(32'sheed9) : $signed(_GEN_15); // @[FFT.scala 34:12]
  assign _GEN_17 = 7'h10 == cnt[6:0] ? $signed(32'shec83) : $signed(_GEN_16); // @[FFT.scala 34:12]
  assign _GEN_18 = 7'h11 == cnt[6:0] ? $signed(32'shea0a) : $signed(_GEN_17); // @[FFT.scala 34:12]
  assign _GEN_19 = 7'h12 == cnt[6:0] ? $signed(32'she76c) : $signed(_GEN_18); // @[FFT.scala 34:12]
  assign _GEN_20 = 7'h13 == cnt[6:0] ? $signed(32'she4aa) : $signed(_GEN_19); // @[FFT.scala 34:12]
  assign _GEN_21 = 7'h14 == cnt[6:0] ? $signed(32'she1c6) : $signed(_GEN_20); // @[FFT.scala 34:12]
  assign _GEN_22 = 7'h15 == cnt[6:0] ? $signed(32'shdebe) : $signed(_GEN_21); // @[FFT.scala 34:12]
  assign _GEN_23 = 7'h16 == cnt[6:0] ? $signed(32'shdb94) : $signed(_GEN_22); // @[FFT.scala 34:12]
  assign _GEN_24 = 7'h17 == cnt[6:0] ? $signed(32'shd848) : $signed(_GEN_23); // @[FFT.scala 34:12]
  assign _GEN_25 = 7'h18 == cnt[6:0] ? $signed(32'shd4db) : $signed(_GEN_24); // @[FFT.scala 34:12]
  assign _GEN_26 = 7'h19 == cnt[6:0] ? $signed(32'shd14d) : $signed(_GEN_25); // @[FFT.scala 34:12]
  assign _GEN_27 = 7'h1a == cnt[6:0] ? $signed(32'shcd9f) : $signed(_GEN_26); // @[FFT.scala 34:12]
  assign _GEN_28 = 7'h1b == cnt[6:0] ? $signed(32'shc9d1) : $signed(_GEN_27); // @[FFT.scala 34:12]
  assign _GEN_29 = 7'h1c == cnt[6:0] ? $signed(32'shc5e4) : $signed(_GEN_28); // @[FFT.scala 34:12]
  assign _GEN_30 = 7'h1d == cnt[6:0] ? $signed(32'shc1d8) : $signed(_GEN_29); // @[FFT.scala 34:12]
  assign _GEN_31 = 7'h1e == cnt[6:0] ? $signed(32'shbdaf) : $signed(_GEN_30); // @[FFT.scala 34:12]
  assign _GEN_32 = 7'h1f == cnt[6:0] ? $signed(32'shb968) : $signed(_GEN_31); // @[FFT.scala 34:12]
  assign _GEN_33 = 7'h20 == cnt[6:0] ? $signed(32'shb505) : $signed(_GEN_32); // @[FFT.scala 34:12]
  assign _GEN_34 = 7'h21 == cnt[6:0] ? $signed(32'shb086) : $signed(_GEN_33); // @[FFT.scala 34:12]
  assign _GEN_35 = 7'h22 == cnt[6:0] ? $signed(32'shabeb) : $signed(_GEN_34); // @[FFT.scala 34:12]
  assign _GEN_36 = 7'h23 == cnt[6:0] ? $signed(32'sha736) : $signed(_GEN_35); // @[FFT.scala 34:12]
  assign _GEN_37 = 7'h24 == cnt[6:0] ? $signed(32'sha268) : $signed(_GEN_36); // @[FFT.scala 34:12]
  assign _GEN_38 = 7'h25 == cnt[6:0] ? $signed(32'sh9d80) : $signed(_GEN_37); // @[FFT.scala 34:12]
  assign _GEN_39 = 7'h26 == cnt[6:0] ? $signed(32'sh9880) : $signed(_GEN_38); // @[FFT.scala 34:12]
  assign _GEN_40 = 7'h27 == cnt[6:0] ? $signed(32'sh9368) : $signed(_GEN_39); // @[FFT.scala 34:12]
  assign _GEN_41 = 7'h28 == cnt[6:0] ? $signed(32'sh8e3a) : $signed(_GEN_40); // @[FFT.scala 34:12]
  assign _GEN_42 = 7'h29 == cnt[6:0] ? $signed(32'sh88f6) : $signed(_GEN_41); // @[FFT.scala 34:12]
  assign _GEN_43 = 7'h2a == cnt[6:0] ? $signed(32'sh839c) : $signed(_GEN_42); // @[FFT.scala 34:12]
  assign _GEN_44 = 7'h2b == cnt[6:0] ? $signed(32'sh7e2f) : $signed(_GEN_43); // @[FFT.scala 34:12]
  assign _GEN_45 = 7'h2c == cnt[6:0] ? $signed(32'sh78ad) : $signed(_GEN_44); // @[FFT.scala 34:12]
  assign _GEN_46 = 7'h2d == cnt[6:0] ? $signed(32'sh731a) : $signed(_GEN_45); // @[FFT.scala 34:12]
  assign _GEN_47 = 7'h2e == cnt[6:0] ? $signed(32'sh6d74) : $signed(_GEN_46); // @[FFT.scala 34:12]
  assign _GEN_48 = 7'h2f == cnt[6:0] ? $signed(32'sh67be) : $signed(_GEN_47); // @[FFT.scala 34:12]
  assign _GEN_49 = 7'h30 == cnt[6:0] ? $signed(32'sh61f8) : $signed(_GEN_48); // @[FFT.scala 34:12]
  assign _GEN_50 = 7'h31 == cnt[6:0] ? $signed(32'sh5c22) : $signed(_GEN_49); // @[FFT.scala 34:12]
  assign _GEN_51 = 7'h32 == cnt[6:0] ? $signed(32'sh563e) : $signed(_GEN_50); // @[FFT.scala 34:12]
  assign _GEN_52 = 7'h33 == cnt[6:0] ? $signed(32'sh504d) : $signed(_GEN_51); // @[FFT.scala 34:12]
  assign _GEN_53 = 7'h34 == cnt[6:0] ? $signed(32'sh4a50) : $signed(_GEN_52); // @[FFT.scala 34:12]
  assign _GEN_54 = 7'h35 == cnt[6:0] ? $signed(32'sh4447) : $signed(_GEN_53); // @[FFT.scala 34:12]
  assign _GEN_55 = 7'h36 == cnt[6:0] ? $signed(32'sh3e34) : $signed(_GEN_54); // @[FFT.scala 34:12]
  assign _GEN_56 = 7'h37 == cnt[6:0] ? $signed(32'sh3817) : $signed(_GEN_55); // @[FFT.scala 34:12]
  assign _GEN_57 = 7'h38 == cnt[6:0] ? $signed(32'sh31f1) : $signed(_GEN_56); // @[FFT.scala 34:12]
  assign _GEN_58 = 7'h39 == cnt[6:0] ? $signed(32'sh2bc4) : $signed(_GEN_57); // @[FFT.scala 34:12]
  assign _GEN_59 = 7'h3a == cnt[6:0] ? $signed(32'sh2590) : $signed(_GEN_58); // @[FFT.scala 34:12]
  assign _GEN_60 = 7'h3b == cnt[6:0] ? $signed(32'sh1f56) : $signed(_GEN_59); // @[FFT.scala 34:12]
  assign _GEN_61 = 7'h3c == cnt[6:0] ? $signed(32'sh1918) : $signed(_GEN_60); // @[FFT.scala 34:12]
  assign _GEN_62 = 7'h3d == cnt[6:0] ? $signed(32'sh12d5) : $signed(_GEN_61); // @[FFT.scala 34:12]
  assign _GEN_63 = 7'h3e == cnt[6:0] ? $signed(32'shc90) : $signed(_GEN_62); // @[FFT.scala 34:12]
  assign _GEN_64 = 7'h3f == cnt[6:0] ? $signed(32'sh648) : $signed(_GEN_63); // @[FFT.scala 34:12]
  assign _GEN_65 = 7'h40 == cnt[6:0] ? $signed(32'sh0) : $signed(_GEN_64); // @[FFT.scala 34:12]
  assign _GEN_66 = 7'h41 == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_65); // @[FFT.scala 34:12]
  assign _GEN_67 = 7'h42 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_66); // @[FFT.scala 34:12]
  assign _GEN_68 = 7'h43 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_67); // @[FFT.scala 34:12]
  assign _GEN_69 = 7'h44 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_68); // @[FFT.scala 34:12]
  assign _GEN_70 = 7'h45 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_69); // @[FFT.scala 34:12]
  assign _GEN_71 = 7'h46 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_70); // @[FFT.scala 34:12]
  assign _GEN_72 = 7'h47 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_71); // @[FFT.scala 34:12]
  assign _GEN_73 = 7'h48 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_72); // @[FFT.scala 34:12]
  assign _GEN_74 = 7'h49 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_73); // @[FFT.scala 34:12]
  assign _GEN_75 = 7'h4a == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_74); // @[FFT.scala 34:12]
  assign _GEN_76 = 7'h4b == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_75); // @[FFT.scala 34:12]
  assign _GEN_77 = 7'h4c == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_76); // @[FFT.scala 34:12]
  assign _GEN_78 = 7'h4d == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_77); // @[FFT.scala 34:12]
  assign _GEN_79 = 7'h4e == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_78); // @[FFT.scala 34:12]
  assign _GEN_80 = 7'h4f == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_79); // @[FFT.scala 34:12]
  assign _GEN_81 = 7'h50 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_80); // @[FFT.scala 34:12]
  assign _GEN_82 = 7'h51 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_81); // @[FFT.scala 34:12]
  assign _GEN_83 = 7'h52 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_82); // @[FFT.scala 34:12]
  assign _GEN_84 = 7'h53 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_83); // @[FFT.scala 34:12]
  assign _GEN_85 = 7'h54 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_84); // @[FFT.scala 34:12]
  assign _GEN_86 = 7'h55 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_85); // @[FFT.scala 34:12]
  assign _GEN_87 = 7'h56 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_86); // @[FFT.scala 34:12]
  assign _GEN_88 = 7'h57 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_87); // @[FFT.scala 34:12]
  assign _GEN_89 = 7'h58 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_88); // @[FFT.scala 34:12]
  assign _GEN_90 = 7'h59 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_89); // @[FFT.scala 34:12]
  assign _GEN_91 = 7'h5a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_90); // @[FFT.scala 34:12]
  assign _GEN_92 = 7'h5b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_91); // @[FFT.scala 34:12]
  assign _GEN_93 = 7'h5c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_92); // @[FFT.scala 34:12]
  assign _GEN_94 = 7'h5d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_93); // @[FFT.scala 34:12]
  assign _GEN_95 = 7'h5e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_94); // @[FFT.scala 34:12]
  assign _GEN_96 = 7'h5f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_95); // @[FFT.scala 34:12]
  assign _GEN_97 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_96); // @[FFT.scala 34:12]
  assign _GEN_98 = 7'h61 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_97); // @[FFT.scala 34:12]
  assign _GEN_99 = 7'h62 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_98); // @[FFT.scala 34:12]
  assign _GEN_100 = 7'h63 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_99); // @[FFT.scala 34:12]
  assign _GEN_101 = 7'h64 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_100); // @[FFT.scala 34:12]
  assign _GEN_102 = 7'h65 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_101); // @[FFT.scala 34:12]
  assign _GEN_103 = 7'h66 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_102); // @[FFT.scala 34:12]
  assign _GEN_104 = 7'h67 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_103); // @[FFT.scala 34:12]
  assign _GEN_105 = 7'h68 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_104); // @[FFT.scala 34:12]
  assign _GEN_106 = 7'h69 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_105); // @[FFT.scala 34:12]
  assign _GEN_107 = 7'h6a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_106); // @[FFT.scala 34:12]
  assign _GEN_108 = 7'h6b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_107); // @[FFT.scala 34:12]
  assign _GEN_109 = 7'h6c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_108); // @[FFT.scala 34:12]
  assign _GEN_110 = 7'h6d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_109); // @[FFT.scala 34:12]
  assign _GEN_111 = 7'h6e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_110); // @[FFT.scala 34:12]
  assign _GEN_112 = 7'h6f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_111); // @[FFT.scala 34:12]
  assign _GEN_113 = 7'h70 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_112); // @[FFT.scala 34:12]
  assign _GEN_114 = 7'h71 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_113); // @[FFT.scala 34:12]
  assign _GEN_115 = 7'h72 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_114); // @[FFT.scala 34:12]
  assign _GEN_116 = 7'h73 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_115); // @[FFT.scala 34:12]
  assign _GEN_117 = 7'h74 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_116); // @[FFT.scala 34:12]
  assign _GEN_118 = 7'h75 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_117); // @[FFT.scala 34:12]
  assign _GEN_119 = 7'h76 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_118); // @[FFT.scala 34:12]
  assign _GEN_120 = 7'h77 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_119); // @[FFT.scala 34:12]
  assign _GEN_121 = 7'h78 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_120); // @[FFT.scala 34:12]
  assign _GEN_122 = 7'h79 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_121); // @[FFT.scala 34:12]
  assign _GEN_123 = 7'h7a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_122); // @[FFT.scala 34:12]
  assign _GEN_124 = 7'h7b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_123); // @[FFT.scala 34:12]
  assign _GEN_125 = 7'h7c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_124); // @[FFT.scala 34:12]
  assign _GEN_126 = 7'h7d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_125); // @[FFT.scala 34:12]
  assign _GEN_127 = 7'h7e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_126); // @[FFT.scala 34:12]
  assign _GEN_130 = 7'h1 == cnt[6:0] ? $signed(-32'sh648) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_131 = 7'h2 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_130); // @[FFT.scala 35:12]
  assign _GEN_132 = 7'h3 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_131); // @[FFT.scala 35:12]
  assign _GEN_133 = 7'h4 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_132); // @[FFT.scala 35:12]
  assign _GEN_134 = 7'h5 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_133); // @[FFT.scala 35:12]
  assign _GEN_135 = 7'h6 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_134); // @[FFT.scala 35:12]
  assign _GEN_136 = 7'h7 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_135); // @[FFT.scala 35:12]
  assign _GEN_137 = 7'h8 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_136); // @[FFT.scala 35:12]
  assign _GEN_138 = 7'h9 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_137); // @[FFT.scala 35:12]
  assign _GEN_139 = 7'ha == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_138); // @[FFT.scala 35:12]
  assign _GEN_140 = 7'hb == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_139); // @[FFT.scala 35:12]
  assign _GEN_141 = 7'hc == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_140); // @[FFT.scala 35:12]
  assign _GEN_142 = 7'hd == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_141); // @[FFT.scala 35:12]
  assign _GEN_143 = 7'he == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_142); // @[FFT.scala 35:12]
  assign _GEN_144 = 7'hf == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_143); // @[FFT.scala 35:12]
  assign _GEN_145 = 7'h10 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_144); // @[FFT.scala 35:12]
  assign _GEN_146 = 7'h11 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_145); // @[FFT.scala 35:12]
  assign _GEN_147 = 7'h12 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_146); // @[FFT.scala 35:12]
  assign _GEN_148 = 7'h13 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_147); // @[FFT.scala 35:12]
  assign _GEN_149 = 7'h14 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_148); // @[FFT.scala 35:12]
  assign _GEN_150 = 7'h15 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_149); // @[FFT.scala 35:12]
  assign _GEN_151 = 7'h16 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_150); // @[FFT.scala 35:12]
  assign _GEN_152 = 7'h17 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_151); // @[FFT.scala 35:12]
  assign _GEN_153 = 7'h18 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_152); // @[FFT.scala 35:12]
  assign _GEN_154 = 7'h19 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_153); // @[FFT.scala 35:12]
  assign _GEN_155 = 7'h1a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_154); // @[FFT.scala 35:12]
  assign _GEN_156 = 7'h1b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_155); // @[FFT.scala 35:12]
  assign _GEN_157 = 7'h1c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_156); // @[FFT.scala 35:12]
  assign _GEN_158 = 7'h1d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_157); // @[FFT.scala 35:12]
  assign _GEN_159 = 7'h1e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_158); // @[FFT.scala 35:12]
  assign _GEN_160 = 7'h1f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_159); // @[FFT.scala 35:12]
  assign _GEN_161 = 7'h20 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_160); // @[FFT.scala 35:12]
  assign _GEN_162 = 7'h21 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_161); // @[FFT.scala 35:12]
  assign _GEN_163 = 7'h22 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_162); // @[FFT.scala 35:12]
  assign _GEN_164 = 7'h23 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_163); // @[FFT.scala 35:12]
  assign _GEN_165 = 7'h24 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_164); // @[FFT.scala 35:12]
  assign _GEN_166 = 7'h25 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_165); // @[FFT.scala 35:12]
  assign _GEN_167 = 7'h26 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_166); // @[FFT.scala 35:12]
  assign _GEN_168 = 7'h27 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_167); // @[FFT.scala 35:12]
  assign _GEN_169 = 7'h28 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_168); // @[FFT.scala 35:12]
  assign _GEN_170 = 7'h29 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_169); // @[FFT.scala 35:12]
  assign _GEN_171 = 7'h2a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_170); // @[FFT.scala 35:12]
  assign _GEN_172 = 7'h2b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_171); // @[FFT.scala 35:12]
  assign _GEN_173 = 7'h2c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_172); // @[FFT.scala 35:12]
  assign _GEN_174 = 7'h2d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_173); // @[FFT.scala 35:12]
  assign _GEN_175 = 7'h2e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_174); // @[FFT.scala 35:12]
  assign _GEN_176 = 7'h2f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_175); // @[FFT.scala 35:12]
  assign _GEN_177 = 7'h30 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_176); // @[FFT.scala 35:12]
  assign _GEN_178 = 7'h31 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_177); // @[FFT.scala 35:12]
  assign _GEN_179 = 7'h32 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_178); // @[FFT.scala 35:12]
  assign _GEN_180 = 7'h33 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_179); // @[FFT.scala 35:12]
  assign _GEN_181 = 7'h34 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_180); // @[FFT.scala 35:12]
  assign _GEN_182 = 7'h35 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_181); // @[FFT.scala 35:12]
  assign _GEN_183 = 7'h36 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_182); // @[FFT.scala 35:12]
  assign _GEN_184 = 7'h37 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_183); // @[FFT.scala 35:12]
  assign _GEN_185 = 7'h38 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_184); // @[FFT.scala 35:12]
  assign _GEN_186 = 7'h39 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_185); // @[FFT.scala 35:12]
  assign _GEN_187 = 7'h3a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_186); // @[FFT.scala 35:12]
  assign _GEN_188 = 7'h3b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_187); // @[FFT.scala 35:12]
  assign _GEN_189 = 7'h3c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_188); // @[FFT.scala 35:12]
  assign _GEN_190 = 7'h3d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_189); // @[FFT.scala 35:12]
  assign _GEN_191 = 7'h3e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_190); // @[FFT.scala 35:12]
  assign _GEN_192 = 7'h3f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_191); // @[FFT.scala 35:12]
  assign _GEN_193 = 7'h40 == cnt[6:0] ? $signed(-32'sh10000) : $signed(_GEN_192); // @[FFT.scala 35:12]
  assign _GEN_194 = 7'h41 == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_193); // @[FFT.scala 35:12]
  assign _GEN_195 = 7'h42 == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_194); // @[FFT.scala 35:12]
  assign _GEN_196 = 7'h43 == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_195); // @[FFT.scala 35:12]
  assign _GEN_197 = 7'h44 == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_196); // @[FFT.scala 35:12]
  assign _GEN_198 = 7'h45 == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_197); // @[FFT.scala 35:12]
  assign _GEN_199 = 7'h46 == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_198); // @[FFT.scala 35:12]
  assign _GEN_200 = 7'h47 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_199); // @[FFT.scala 35:12]
  assign _GEN_201 = 7'h48 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_200); // @[FFT.scala 35:12]
  assign _GEN_202 = 7'h49 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_201); // @[FFT.scala 35:12]
  assign _GEN_203 = 7'h4a == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_202); // @[FFT.scala 35:12]
  assign _GEN_204 = 7'h4b == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_203); // @[FFT.scala 35:12]
  assign _GEN_205 = 7'h4c == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_204); // @[FFT.scala 35:12]
  assign _GEN_206 = 7'h4d == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_205); // @[FFT.scala 35:12]
  assign _GEN_207 = 7'h4e == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_206); // @[FFT.scala 35:12]
  assign _GEN_208 = 7'h4f == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_207); // @[FFT.scala 35:12]
  assign _GEN_209 = 7'h50 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_208); // @[FFT.scala 35:12]
  assign _GEN_210 = 7'h51 == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_209); // @[FFT.scala 35:12]
  assign _GEN_211 = 7'h52 == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_210); // @[FFT.scala 35:12]
  assign _GEN_212 = 7'h53 == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_211); // @[FFT.scala 35:12]
  assign _GEN_213 = 7'h54 == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_212); // @[FFT.scala 35:12]
  assign _GEN_214 = 7'h55 == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_213); // @[FFT.scala 35:12]
  assign _GEN_215 = 7'h56 == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_214); // @[FFT.scala 35:12]
  assign _GEN_216 = 7'h57 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_215); // @[FFT.scala 35:12]
  assign _GEN_217 = 7'h58 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_216); // @[FFT.scala 35:12]
  assign _GEN_218 = 7'h59 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_217); // @[FFT.scala 35:12]
  assign _GEN_219 = 7'h5a == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_218); // @[FFT.scala 35:12]
  assign _GEN_220 = 7'h5b == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_219); // @[FFT.scala 35:12]
  assign _GEN_221 = 7'h5c == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_220); // @[FFT.scala 35:12]
  assign _GEN_222 = 7'h5d == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_221); // @[FFT.scala 35:12]
  assign _GEN_223 = 7'h5e == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_222); // @[FFT.scala 35:12]
  assign _GEN_224 = 7'h5f == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_223); // @[FFT.scala 35:12]
  assign _GEN_225 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_224); // @[FFT.scala 35:12]
  assign _GEN_226 = 7'h61 == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_225); // @[FFT.scala 35:12]
  assign _GEN_227 = 7'h62 == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_226); // @[FFT.scala 35:12]
  assign _GEN_228 = 7'h63 == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_227); // @[FFT.scala 35:12]
  assign _GEN_229 = 7'h64 == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_228); // @[FFT.scala 35:12]
  assign _GEN_230 = 7'h65 == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_229); // @[FFT.scala 35:12]
  assign _GEN_231 = 7'h66 == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_230); // @[FFT.scala 35:12]
  assign _GEN_232 = 7'h67 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_231); // @[FFT.scala 35:12]
  assign _GEN_233 = 7'h68 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_232); // @[FFT.scala 35:12]
  assign _GEN_234 = 7'h69 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_233); // @[FFT.scala 35:12]
  assign _GEN_235 = 7'h6a == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_234); // @[FFT.scala 35:12]
  assign _GEN_236 = 7'h6b == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_235); // @[FFT.scala 35:12]
  assign _GEN_237 = 7'h6c == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_236); // @[FFT.scala 35:12]
  assign _GEN_238 = 7'h6d == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_237); // @[FFT.scala 35:12]
  assign _GEN_239 = 7'h6e == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_238); // @[FFT.scala 35:12]
  assign _GEN_240 = 7'h6f == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_239); // @[FFT.scala 35:12]
  assign _GEN_241 = 7'h70 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_240); // @[FFT.scala 35:12]
  assign _GEN_242 = 7'h71 == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_241); // @[FFT.scala 35:12]
  assign _GEN_243 = 7'h72 == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_242); // @[FFT.scala 35:12]
  assign _GEN_244 = 7'h73 == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_243); // @[FFT.scala 35:12]
  assign _GEN_245 = 7'h74 == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_244); // @[FFT.scala 35:12]
  assign _GEN_246 = 7'h75 == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_245); // @[FFT.scala 35:12]
  assign _GEN_247 = 7'h76 == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_246); // @[FFT.scala 35:12]
  assign _GEN_248 = 7'h77 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_247); // @[FFT.scala 35:12]
  assign _GEN_249 = 7'h78 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_248); // @[FFT.scala 35:12]
  assign _GEN_250 = 7'h79 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_249); // @[FFT.scala 35:12]
  assign _GEN_251 = 7'h7a == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_250); // @[FFT.scala 35:12]
  assign _GEN_252 = 7'h7b == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_251); // @[FFT.scala 35:12]
  assign _GEN_253 = 7'h7c == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_252); // @[FFT.scala 35:12]
  assign _GEN_254 = 7'h7d == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_253); // @[FFT.scala 35:12]
  assign _GEN_255 = 7'h7e == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_254); // @[FFT.scala 35:12]
  assign _GEN_642 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_643 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_642); // @[FFT.scala 34:12]
  assign _GEN_644 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_643); // @[FFT.scala 34:12]
  assign _GEN_645 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_644); // @[FFT.scala 34:12]
  assign _GEN_646 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_645); // @[FFT.scala 34:12]
  assign _GEN_647 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_646); // @[FFT.scala 34:12]
  assign _GEN_648 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_647); // @[FFT.scala 34:12]
  assign _GEN_649 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_648); // @[FFT.scala 34:12]
  assign _GEN_650 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_649); // @[FFT.scala 34:12]
  assign _GEN_651 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_650); // @[FFT.scala 34:12]
  assign _GEN_652 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_651); // @[FFT.scala 34:12]
  assign _GEN_653 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_652); // @[FFT.scala 34:12]
  assign _GEN_654 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_653); // @[FFT.scala 34:12]
  assign _GEN_655 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_654); // @[FFT.scala 34:12]
  assign _GEN_656 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_655); // @[FFT.scala 34:12]
  assign _GEN_657 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_656); // @[FFT.scala 34:12]
  assign _GEN_658 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_657); // @[FFT.scala 34:12]
  assign _GEN_659 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_658); // @[FFT.scala 34:12]
  assign _GEN_660 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_659); // @[FFT.scala 34:12]
  assign _GEN_661 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_660); // @[FFT.scala 34:12]
  assign _GEN_662 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_661); // @[FFT.scala 34:12]
  assign _GEN_663 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_662); // @[FFT.scala 34:12]
  assign _GEN_664 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_663); // @[FFT.scala 34:12]
  assign _GEN_665 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_664); // @[FFT.scala 34:12]
  assign _GEN_666 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_665); // @[FFT.scala 34:12]
  assign _GEN_667 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_666); // @[FFT.scala 34:12]
  assign _GEN_668 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_667); // @[FFT.scala 34:12]
  assign _GEN_669 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_668); // @[FFT.scala 34:12]
  assign _GEN_670 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_669); // @[FFT.scala 34:12]
  assign _GEN_671 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_670); // @[FFT.scala 34:12]
  assign _GEN_672 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_671); // @[FFT.scala 34:12]
  assign _GEN_673 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_672); // @[FFT.scala 34:12]
  assign _GEN_674 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_673); // @[FFT.scala 34:12]
  assign _GEN_675 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_674); // @[FFT.scala 34:12]
  assign _GEN_676 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_675); // @[FFT.scala 34:12]
  assign _GEN_677 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_676); // @[FFT.scala 34:12]
  assign _GEN_678 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_677); // @[FFT.scala 34:12]
  assign _GEN_679 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_678); // @[FFT.scala 34:12]
  assign _GEN_680 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_679); // @[FFT.scala 34:12]
  assign _GEN_681 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_680); // @[FFT.scala 34:12]
  assign _GEN_682 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_681); // @[FFT.scala 34:12]
  assign _GEN_683 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_682); // @[FFT.scala 34:12]
  assign _GEN_684 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_683); // @[FFT.scala 34:12]
  assign _GEN_685 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_684); // @[FFT.scala 34:12]
  assign _GEN_686 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_685); // @[FFT.scala 34:12]
  assign _GEN_687 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_686); // @[FFT.scala 34:12]
  assign _GEN_688 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_687); // @[FFT.scala 34:12]
  assign _GEN_689 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_688); // @[FFT.scala 34:12]
  assign _GEN_690 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_689); // @[FFT.scala 34:12]
  assign _GEN_691 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_690); // @[FFT.scala 34:12]
  assign _GEN_692 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_691); // @[FFT.scala 34:12]
  assign _GEN_693 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_692); // @[FFT.scala 34:12]
  assign _GEN_694 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_693); // @[FFT.scala 34:12]
  assign _GEN_695 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_694); // @[FFT.scala 34:12]
  assign _GEN_696 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_695); // @[FFT.scala 34:12]
  assign _GEN_697 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_696); // @[FFT.scala 34:12]
  assign _GEN_698 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_697); // @[FFT.scala 34:12]
  assign _GEN_699 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_698); // @[FFT.scala 34:12]
  assign _GEN_700 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_699); // @[FFT.scala 34:12]
  assign _GEN_701 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_700); // @[FFT.scala 34:12]
  assign _GEN_702 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_701); // @[FFT.scala 34:12]
  assign _GEN_703 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_702); // @[FFT.scala 34:12]
  assign _GEN_706 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_707 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_706); // @[FFT.scala 35:12]
  assign _GEN_708 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_707); // @[FFT.scala 35:12]
  assign _GEN_709 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_708); // @[FFT.scala 35:12]
  assign _GEN_710 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_709); // @[FFT.scala 35:12]
  assign _GEN_711 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_710); // @[FFT.scala 35:12]
  assign _GEN_712 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_711); // @[FFT.scala 35:12]
  assign _GEN_713 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_712); // @[FFT.scala 35:12]
  assign _GEN_714 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_713); // @[FFT.scala 35:12]
  assign _GEN_715 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_714); // @[FFT.scala 35:12]
  assign _GEN_716 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_715); // @[FFT.scala 35:12]
  assign _GEN_717 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_716); // @[FFT.scala 35:12]
  assign _GEN_718 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_717); // @[FFT.scala 35:12]
  assign _GEN_719 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_718); // @[FFT.scala 35:12]
  assign _GEN_720 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_719); // @[FFT.scala 35:12]
  assign _GEN_721 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_720); // @[FFT.scala 35:12]
  assign _GEN_722 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_721); // @[FFT.scala 35:12]
  assign _GEN_723 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_722); // @[FFT.scala 35:12]
  assign _GEN_724 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_723); // @[FFT.scala 35:12]
  assign _GEN_725 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_724); // @[FFT.scala 35:12]
  assign _GEN_726 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_725); // @[FFT.scala 35:12]
  assign _GEN_727 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_726); // @[FFT.scala 35:12]
  assign _GEN_728 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_727); // @[FFT.scala 35:12]
  assign _GEN_729 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_728); // @[FFT.scala 35:12]
  assign _GEN_730 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_729); // @[FFT.scala 35:12]
  assign _GEN_731 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_730); // @[FFT.scala 35:12]
  assign _GEN_732 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_731); // @[FFT.scala 35:12]
  assign _GEN_733 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_732); // @[FFT.scala 35:12]
  assign _GEN_734 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_733); // @[FFT.scala 35:12]
  assign _GEN_735 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_734); // @[FFT.scala 35:12]
  assign _GEN_736 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_735); // @[FFT.scala 35:12]
  assign _GEN_737 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_736); // @[FFT.scala 35:12]
  assign _GEN_738 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_737); // @[FFT.scala 35:12]
  assign _GEN_739 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_738); // @[FFT.scala 35:12]
  assign _GEN_740 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_739); // @[FFT.scala 35:12]
  assign _GEN_741 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_740); // @[FFT.scala 35:12]
  assign _GEN_742 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_741); // @[FFT.scala 35:12]
  assign _GEN_743 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_742); // @[FFT.scala 35:12]
  assign _GEN_744 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_743); // @[FFT.scala 35:12]
  assign _GEN_745 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_744); // @[FFT.scala 35:12]
  assign _GEN_746 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_745); // @[FFT.scala 35:12]
  assign _GEN_747 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_746); // @[FFT.scala 35:12]
  assign _GEN_748 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_747); // @[FFT.scala 35:12]
  assign _GEN_749 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_748); // @[FFT.scala 35:12]
  assign _GEN_750 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_749); // @[FFT.scala 35:12]
  assign _GEN_751 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_750); // @[FFT.scala 35:12]
  assign _GEN_752 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_751); // @[FFT.scala 35:12]
  assign _GEN_753 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_752); // @[FFT.scala 35:12]
  assign _GEN_754 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_753); // @[FFT.scala 35:12]
  assign _GEN_755 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_754); // @[FFT.scala 35:12]
  assign _GEN_756 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_755); // @[FFT.scala 35:12]
  assign _GEN_757 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_756); // @[FFT.scala 35:12]
  assign _GEN_758 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_757); // @[FFT.scala 35:12]
  assign _GEN_759 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_758); // @[FFT.scala 35:12]
  assign _GEN_760 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_759); // @[FFT.scala 35:12]
  assign _GEN_761 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_760); // @[FFT.scala 35:12]
  assign _GEN_762 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_761); // @[FFT.scala 35:12]
  assign _GEN_763 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_762); // @[FFT.scala 35:12]
  assign _GEN_764 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_763); // @[FFT.scala 35:12]
  assign _GEN_765 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_764); // @[FFT.scala 35:12]
  assign _GEN_766 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_765); // @[FFT.scala 35:12]
  assign _GEN_767 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_766); // @[FFT.scala 35:12]
  assign _GEN_962 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_963 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_962); // @[FFT.scala 34:12]
  assign _GEN_964 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_963); // @[FFT.scala 34:12]
  assign _GEN_965 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_964); // @[FFT.scala 34:12]
  assign _GEN_966 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_965); // @[FFT.scala 34:12]
  assign _GEN_967 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_966); // @[FFT.scala 34:12]
  assign _GEN_968 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_967); // @[FFT.scala 34:12]
  assign _GEN_969 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_968); // @[FFT.scala 34:12]
  assign _GEN_970 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_969); // @[FFT.scala 34:12]
  assign _GEN_971 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_970); // @[FFT.scala 34:12]
  assign _GEN_972 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_971); // @[FFT.scala 34:12]
  assign _GEN_973 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_972); // @[FFT.scala 34:12]
  assign _GEN_974 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_973); // @[FFT.scala 34:12]
  assign _GEN_975 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_974); // @[FFT.scala 34:12]
  assign _GEN_976 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_975); // @[FFT.scala 34:12]
  assign _GEN_977 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_976); // @[FFT.scala 34:12]
  assign _GEN_978 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_977); // @[FFT.scala 34:12]
  assign _GEN_979 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_978); // @[FFT.scala 34:12]
  assign _GEN_980 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_979); // @[FFT.scala 34:12]
  assign _GEN_981 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_980); // @[FFT.scala 34:12]
  assign _GEN_982 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_981); // @[FFT.scala 34:12]
  assign _GEN_983 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_982); // @[FFT.scala 34:12]
  assign _GEN_984 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_983); // @[FFT.scala 34:12]
  assign _GEN_985 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_984); // @[FFT.scala 34:12]
  assign _GEN_986 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_985); // @[FFT.scala 34:12]
  assign _GEN_987 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_986); // @[FFT.scala 34:12]
  assign _GEN_988 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_987); // @[FFT.scala 34:12]
  assign _GEN_989 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_988); // @[FFT.scala 34:12]
  assign _GEN_990 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_989); // @[FFT.scala 34:12]
  assign _GEN_991 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_990); // @[FFT.scala 34:12]
  assign _GEN_994 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_995 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_994); // @[FFT.scala 35:12]
  assign _GEN_996 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_995); // @[FFT.scala 35:12]
  assign _GEN_997 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_996); // @[FFT.scala 35:12]
  assign _GEN_998 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_997); // @[FFT.scala 35:12]
  assign _GEN_999 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_998); // @[FFT.scala 35:12]
  assign _GEN_1000 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_999); // @[FFT.scala 35:12]
  assign _GEN_1001 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_1000); // @[FFT.scala 35:12]
  assign _GEN_1002 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_1001); // @[FFT.scala 35:12]
  assign _GEN_1003 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_1002); // @[FFT.scala 35:12]
  assign _GEN_1004 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_1003); // @[FFT.scala 35:12]
  assign _GEN_1005 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_1004); // @[FFT.scala 35:12]
  assign _GEN_1006 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_1005); // @[FFT.scala 35:12]
  assign _GEN_1007 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_1006); // @[FFT.scala 35:12]
  assign _GEN_1008 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_1007); // @[FFT.scala 35:12]
  assign _GEN_1009 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_1008); // @[FFT.scala 35:12]
  assign _GEN_1010 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_1009); // @[FFT.scala 35:12]
  assign _GEN_1011 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_1010); // @[FFT.scala 35:12]
  assign _GEN_1012 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_1011); // @[FFT.scala 35:12]
  assign _GEN_1013 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_1012); // @[FFT.scala 35:12]
  assign _GEN_1014 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_1013); // @[FFT.scala 35:12]
  assign _GEN_1015 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_1014); // @[FFT.scala 35:12]
  assign _GEN_1016 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_1015); // @[FFT.scala 35:12]
  assign _GEN_1017 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_1016); // @[FFT.scala 35:12]
  assign _GEN_1018 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_1017); // @[FFT.scala 35:12]
  assign _GEN_1019 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1018); // @[FFT.scala 35:12]
  assign _GEN_1020 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_1019); // @[FFT.scala 35:12]
  assign _GEN_1021 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_1020); // @[FFT.scala 35:12]
  assign _GEN_1022 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_1021); // @[FFT.scala 35:12]
  assign _GEN_1023 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_1022); // @[FFT.scala 35:12]
  assign _GEN_1122 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1123 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_1122); // @[FFT.scala 34:12]
  assign _GEN_1124 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_1123); // @[FFT.scala 34:12]
  assign _GEN_1125 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_1124); // @[FFT.scala 34:12]
  assign _GEN_1126 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_1125); // @[FFT.scala 34:12]
  assign _GEN_1127 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_1126); // @[FFT.scala 34:12]
  assign _GEN_1128 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_1127); // @[FFT.scala 34:12]
  assign _GEN_1129 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_1128); // @[FFT.scala 34:12]
  assign _GEN_1130 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_1129); // @[FFT.scala 34:12]
  assign _GEN_1131 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_1130); // @[FFT.scala 34:12]
  assign _GEN_1132 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1131); // @[FFT.scala 34:12]
  assign _GEN_1133 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_1132); // @[FFT.scala 34:12]
  assign _GEN_1134 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_1133); // @[FFT.scala 34:12]
  assign _GEN_1135 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_1134); // @[FFT.scala 34:12]
  assign _GEN_1138 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1139 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_1138); // @[FFT.scala 35:12]
  assign _GEN_1140 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1139); // @[FFT.scala 35:12]
  assign _GEN_1141 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_1140); // @[FFT.scala 35:12]
  assign _GEN_1142 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_1141); // @[FFT.scala 35:12]
  assign _GEN_1143 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_1142); // @[FFT.scala 35:12]
  assign _GEN_1144 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_1143); // @[FFT.scala 35:12]
  assign _GEN_1145 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_1144); // @[FFT.scala 35:12]
  assign _GEN_1146 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_1145); // @[FFT.scala 35:12]
  assign _GEN_1147 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_1146); // @[FFT.scala 35:12]
  assign _GEN_1148 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_1147); // @[FFT.scala 35:12]
  assign _GEN_1149 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_1148); // @[FFT.scala 35:12]
  assign _GEN_1150 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1149); // @[FFT.scala 35:12]
  assign _GEN_1151 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_1150); // @[FFT.scala 35:12]
  assign _GEN_1202 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1203 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_1202); // @[FFT.scala 34:12]
  assign _GEN_1204 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_1203); // @[FFT.scala 34:12]
  assign _GEN_1205 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_1204); // @[FFT.scala 34:12]
  assign _GEN_1206 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_1205); // @[FFT.scala 34:12]
  assign _GEN_1207 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_1206); // @[FFT.scala 34:12]
  assign _GEN_1210 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1211 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_1210); // @[FFT.scala 35:12]
  assign _GEN_1212 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_1211); // @[FFT.scala 35:12]
  assign _GEN_1213 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_1212); // @[FFT.scala 35:12]
  assign _GEN_1214 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_1213); // @[FFT.scala 35:12]
  assign _GEN_1215 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_1214); // @[FFT.scala 35:12]
  assign _GEN_1242 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1243 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_1242); // @[FFT.scala 34:12]
  assign _GEN_1246 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1247 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_1246); // @[FFT.scala 35:12]
  assign io_dOut1_re = _T_544_re; // @[FFT.scala 62:12]
  assign io_dOut1_im = _T_544_im; // @[FFT.scala 62:12]
  assign io_dOut2_re = _T_545_re; // @[FFT.scala 63:12]
  assign io_dOut2_im = _T_545_im; // @[FFT.scala 63:12]
  assign io_dout_valid = _T_801; // @[FFT.scala 64:17]
  assign Butterfly_io_in1_re = _T_259_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_259_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = io_dIn_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = 7'h7f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_127); // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = 7'h7f == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_255); // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_324_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_324_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cnt[6]; // @[Butterfly.scala 113:17]
  assign Butterfly_1_io_in1_re = _T_392_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_392_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_703); // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_767); // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_425_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_425_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cnt[5]; // @[Butterfly.scala 113:17]
  assign Butterfly_2_io_in1_re = _T_461_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_461_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_991); // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_1023); // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_478_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_478_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cnt[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_3_io_in1_re = _T_498_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_498_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_1135); // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_1151); // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_507_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_507_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cnt[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_519_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_519_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_1207); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_1215); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_524_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_524_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cnt[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_532_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_532_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_1243); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_1247); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_535_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_535_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cnt[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_541_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_541_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_543_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_543_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cnt[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_6_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_6_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_6_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_6_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_132_re = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_132_im = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_133_re = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_133_im = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_134_re = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_134_im = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_135_re = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_135_im = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_136_re = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_136_im = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_137_re = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_137_im = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_138_re = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_138_im = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_139_re = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_139_im = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_140_re = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_140_im = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_141_re = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_141_im = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_142_re = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_142_im = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_143_re = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_143_im = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_144_re = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_144_im = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_145_re = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_145_im = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_146_re = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_146_im = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_147_re = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_147_im = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_148_re = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_148_im = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_149_re = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_149_im = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_150_re = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_150_im = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_151_re = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_151_im = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_152_re = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_152_im = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_153_re = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_153_im = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_154_re = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_154_im = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_155_re = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_155_im = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_156_re = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_156_im = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_157_re = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_157_im = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_158_re = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_158_im = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_159_re = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_159_im = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_160_re = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_160_im = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_161_re = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_161_im = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_162_re = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_162_im = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_163_re = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_163_im = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_164_re = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_164_im = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_165_re = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_165_im = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_166_re = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_166_im = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_167_re = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_167_im = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_168_re = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_168_im = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_169_re = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_169_im = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_170_re = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_170_im = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_171_re = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_171_im = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_172_re = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_172_im = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_173_re = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_173_im = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_174_re = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_174_im = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_175_re = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_175_im = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_176_re = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_176_im = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_177_re = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_177_im = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_178_re = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_178_im = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_179_re = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_179_im = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_180_re = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_180_im = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_181_re = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_181_im = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_182_re = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_182_im = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_183_re = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_183_im = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_184_re = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_184_im = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_185_re = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_185_im = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_186_re = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_186_im = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_187_re = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_187_im = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_188_re = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_188_im = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_189_re = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_189_im = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_190_re = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_190_im = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_191_re = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_191_im = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_192_re = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_192_im = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_193_re = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_193_im = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_194_re = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_194_im = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_195_re = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_195_im = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_196_re = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_196_im = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_197_re = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_197_im = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_198_re = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_198_im = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_199_re = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_199_im = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_200_re = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_200_im = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_201_re = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_201_im = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_202_re = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_202_im = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_203_re = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_203_im = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_204_re = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_204_im = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_205_re = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_205_im = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_206_re = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_206_im = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_207_re = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_207_im = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_208_re = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_208_im = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_209_re = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_209_im = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_210_re = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_210_im = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_211_re = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_211_im = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_212_re = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_212_im = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_213_re = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_213_im = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_214_re = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_214_im = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_215_re = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_215_im = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_216_re = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_216_im = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_217_re = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_217_im = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_218_re = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_218_im = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_219_re = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_219_im = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_220_re = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_220_im = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_221_re = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_221_im = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_222_re = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_222_im = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_223_re = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_223_im = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_224_re = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_224_im = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_225_re = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_225_im = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_226_re = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_226_im = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_227_re = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_227_im = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_228_re = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_228_im = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_229_re = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_229_im = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_230_re = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_230_im = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_231_re = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_231_im = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_232_re = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_232_im = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_233_re = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_233_im = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_234_re = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_234_im = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_235_re = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_235_im = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_236_re = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_236_im = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_237_re = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_237_im = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_238_re = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_238_im = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_239_re = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_239_im = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_240_re = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_240_im = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_241_re = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_241_im = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_242_re = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_242_im = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_243_re = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_243_im = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_244_re = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_244_im = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_245_re = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_245_im = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_246_re = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_246_im = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_247_re = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_247_im = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_248_re = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_248_im = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_249_re = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_249_im = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_250_re = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_250_im = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_251_re = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_251_im = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_252_re = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_252_im = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_253_re = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_253_im = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_254_re = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_254_im = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_255_re = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_255_im = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_256_re = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_256_im = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_257_re = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_257_im = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_258_re = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_258_im = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_259_re = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_259_im = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_261_re = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_261_im = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_262_re = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_262_im = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_263_re = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_263_im = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_264_re = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_264_im = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_265_re = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_265_im = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_266_re = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_266_im = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_267_re = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_267_im = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_268_re = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_268_im = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_269_re = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_269_im = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_270_re = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_270_im = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_271_re = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_271_im = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_272_re = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_272_im = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_273_re = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_273_im = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_274_re = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_274_im = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_275_re = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_275_im = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_276_re = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_276_im = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_277_re = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_277_im = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_278_re = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_278_im = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_279_re = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_279_im = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_280_re = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_280_im = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_281_re = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_281_im = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_282_re = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_282_im = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_283_re = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_283_im = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_284_re = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_284_im = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_285_re = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_285_im = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_286_re = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_286_im = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_287_re = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_287_im = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_288_re = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_288_im = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_289_re = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_289_im = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_290_re = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_290_im = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_291_re = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_291_im = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_292_re = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_292_im = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_293_re = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_293_im = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_294_re = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_294_im = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_295_re = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_295_im = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_296_re = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_296_im = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_297_re = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_297_im = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_298_re = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_298_im = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_299_re = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_299_im = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_300_re = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_300_im = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_301_re = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_301_im = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_302_re = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_302_im = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_303_re = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_303_im = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_304_re = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_304_im = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_305_re = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_305_im = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_306_re = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_306_im = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_307_re = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_307_im = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_308_re = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_308_im = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_309_re = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_309_im = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_310_re = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_310_im = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_311_re = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_311_im = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_312_re = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_312_im = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_313_re = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_313_im = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_314_re = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_314_im = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_315_re = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_315_im = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_316_re = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_316_im = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_317_re = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_317_im = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_318_re = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_318_im = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_319_re = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_319_im = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_320_re = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_320_im = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_321_re = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_321_im = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_322_re = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_322_im = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_323_re = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_323_im = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_324_re = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_324_im = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_329_re = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_329_im = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_330_re = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_330_im = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_331_re = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_331_im = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_332_re = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_332_im = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_333_re = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_333_im = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_334_re = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_334_im = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_335_re = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_335_im = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_336_re = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_336_im = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_337_re = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_337_im = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_338_re = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_338_im = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_339_re = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_339_im = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_340_re = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_340_im = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_341_re = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_341_im = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_342_re = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_342_im = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_343_re = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_343_im = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_344_re = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_344_im = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_345_re = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_345_im = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_346_re = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_346_im = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_347_re = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_347_im = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_348_re = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_348_im = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_349_re = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_349_im = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_350_re = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_350_im = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_351_re = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_351_im = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_352_re = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_352_im = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_353_re = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_353_im = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_354_re = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_354_im = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_355_re = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_355_im = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_356_re = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_356_im = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_357_re = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_357_im = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_358_re = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_358_im = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_359_re = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_359_im = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_360_re = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_360_im = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_361_re = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_361_im = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_362_re = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_362_im = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_363_re = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_363_im = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_364_re = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_364_im = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_365_re = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_365_im = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_366_re = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_366_im = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_367_re = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_367_im = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_368_re = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_368_im = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_369_re = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_369_im = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_370_re = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_370_im = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_371_re = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_371_im = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_372_re = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_372_im = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_373_re = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_373_im = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_374_re = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_374_im = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_375_re = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_375_im = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_376_re = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_376_im = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_377_re = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_377_im = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_378_re = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_378_im = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_379_re = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_379_im = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_380_re = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_380_im = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_381_re = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_381_im = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_382_re = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_382_im = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_383_re = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_383_im = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_384_re = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_384_im = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_385_re = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_385_im = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_386_re = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_386_im = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_387_re = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_387_im = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_388_re = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_388_im = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_389_re = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_389_im = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_390_re = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_390_im = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_391_re = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_391_im = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_392_re = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_392_im = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_394_re = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_394_im = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_395_re = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_395_im = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_396_re = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_396_im = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_397_re = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_397_im = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_398_re = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_398_im = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_399_re = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_399_im = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_400_re = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_400_im = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_401_re = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_401_im = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_402_re = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_402_im = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_403_re = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_403_im = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_404_re = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_404_im = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_405_re = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_405_im = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_406_re = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_406_im = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_407_re = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_407_im = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_408_re = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_408_im = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_409_re = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_409_im = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_410_re = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_410_im = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_411_re = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_411_im = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_412_re = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_412_im = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_413_re = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_413_im = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_414_re = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_414_im = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_415_re = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_415_im = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_416_re = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_416_im = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_417_re = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_417_im = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_418_re = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_418_im = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_419_re = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_419_im = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_420_re = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_420_im = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_421_re = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_421_im = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_422_re = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_422_im = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_423_re = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_423_im = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_424_re = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_424_im = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_425_re = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_425_im = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_430_re = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_430_im = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_431_re = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_431_im = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_432_re = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_432_im = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_433_re = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_433_im = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_434_re = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_434_im = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_435_re = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_435_im = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_436_re = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_436_im = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_437_re = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_437_im = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_438_re = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_438_im = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_439_re = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_439_im = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_440_re = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_440_im = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_441_re = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_441_im = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_442_re = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_442_im = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_443_re = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_443_im = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_444_re = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_444_im = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_445_re = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_445_im = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_446_re = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_446_im = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_447_re = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_447_im = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_448_re = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_448_im = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_449_re = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_449_im = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_450_re = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_450_im = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_451_re = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_451_im = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_452_re = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_452_im = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_453_re = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_453_im = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_454_re = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_454_im = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_455_re = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_455_im = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_456_re = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_456_im = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_457_re = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_457_im = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_458_re = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_458_im = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_459_re = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_459_im = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_460_re = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_460_im = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_461_re = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_461_im = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_463_re = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_463_im = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_464_re = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_464_im = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_465_re = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_465_im = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_466_re = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_466_im = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_467_re = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_467_im = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_468_re = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_468_im = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_469_re = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_469_im = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_470_re = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_470_im = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_471_re = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_471_im = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_472_re = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_472_im = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_473_re = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_473_im = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_474_re = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_474_im = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_475_re = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_475_im = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_476_re = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_476_im = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_477_re = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_477_im = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_478_re = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_478_im = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_483_re = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_483_im = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_484_re = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_484_im = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_485_re = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_485_im = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_486_re = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_486_im = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_487_re = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_487_im = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_488_re = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_488_im = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_489_re = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_489_im = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_490_re = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_490_im = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_491_re = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_491_im = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_492_re = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_492_im = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_493_re = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_493_im = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_494_re = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_494_im = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_495_re = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_495_im = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_496_re = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_496_im = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_497_re = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_497_im = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_498_re = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_498_im = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_500_re = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_500_im = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_501_re = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_501_im = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_502_re = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_502_im = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_503_re = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_503_im = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_504_re = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_504_im = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_505_re = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_505_im = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_506_re = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_506_im = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_507_re = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_507_im = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_512_re = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_512_im = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_513_re = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_513_im = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_514_re = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_514_im = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_515_re = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_515_im = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_516_re = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_516_im = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_517_re = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_517_im = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_518_re = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_518_im = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_519_re = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_519_im = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_521_re = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_521_im = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_522_re = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_522_im = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_523_re = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_523_im = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_524_re = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_524_im = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_529_re = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_529_im = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_530_re = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_530_im = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_531_re = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_531_im = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_532_re = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_532_im = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_534_re = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_534_im = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_535_re = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_535_im = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_540_re = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_540_im = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_541_re = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_541_im = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_543_re = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_543_im = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  out1D1_re = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  out1D1_im = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_544_re = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_544_im = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_545_re = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_545_im = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_546 = _RAND_769[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_547 = _RAND_770[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_548 = _RAND_771[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_549 = _RAND_772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_550 = _RAND_773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_551 = _RAND_774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_552 = _RAND_775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_553 = _RAND_776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_554 = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_555 = _RAND_778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_556 = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_557 = _RAND_780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_558 = _RAND_781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_559 = _RAND_782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_560 = _RAND_783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_561 = _RAND_784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_562 = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_563 = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_564 = _RAND_787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_565 = _RAND_788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_566 = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_567 = _RAND_790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_568 = _RAND_791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_569 = _RAND_792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_570 = _RAND_793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_571 = _RAND_794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_572 = _RAND_795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_573 = _RAND_796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_574 = _RAND_797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_575 = _RAND_798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_576 = _RAND_799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_577 = _RAND_800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_578 = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_579 = _RAND_802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_580 = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_581 = _RAND_804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_582 = _RAND_805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_583 = _RAND_806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_584 = _RAND_807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_585 = _RAND_808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_586 = _RAND_809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_587 = _RAND_810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_588 = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_589 = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_590 = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_591 = _RAND_814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_592 = _RAND_815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_593 = _RAND_816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_594 = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_595 = _RAND_818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_596 = _RAND_819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_597 = _RAND_820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_598 = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_599 = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_600 = _RAND_823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_601 = _RAND_824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_602 = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_603 = _RAND_826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_604 = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_605 = _RAND_828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_606 = _RAND_829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_607 = _RAND_830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_608 = _RAND_831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_609 = _RAND_832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_610 = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_611 = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_612 = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_613 = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_614 = _RAND_837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_615 = _RAND_838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_616 = _RAND_839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_617 = _RAND_840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_618 = _RAND_841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_619 = _RAND_842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_620 = _RAND_843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_621 = _RAND_844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_622 = _RAND_845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_623 = _RAND_846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_624 = _RAND_847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_625 = _RAND_848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_626 = _RAND_849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_627 = _RAND_850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_628 = _RAND_851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_629 = _RAND_852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_630 = _RAND_853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_631 = _RAND_854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_632 = _RAND_855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_633 = _RAND_856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_634 = _RAND_857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_635 = _RAND_858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_636 = _RAND_859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_637 = _RAND_860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_638 = _RAND_861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_639 = _RAND_862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_640 = _RAND_863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_641 = _RAND_864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_642 = _RAND_865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_643 = _RAND_866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_644 = _RAND_867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_645 = _RAND_868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_646 = _RAND_869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_647 = _RAND_870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_648 = _RAND_871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_649 = _RAND_872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_650 = _RAND_873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_651 = _RAND_874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_652 = _RAND_875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_653 = _RAND_876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_654 = _RAND_877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_655 = _RAND_878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_656 = _RAND_879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_657 = _RAND_880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_658 = _RAND_881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_659 = _RAND_882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_660 = _RAND_883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_661 = _RAND_884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_662 = _RAND_885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_663 = _RAND_886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_664 = _RAND_887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_665 = _RAND_888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_666 = _RAND_889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_667 = _RAND_890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_668 = _RAND_891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_669 = _RAND_892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_670 = _RAND_893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_671 = _RAND_894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_672 = _RAND_895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_673 = _RAND_896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_674 = _RAND_897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_675 = _RAND_898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_676 = _RAND_899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_677 = _RAND_900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_678 = _RAND_901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_679 = _RAND_902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_680 = _RAND_903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_681 = _RAND_904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_682 = _RAND_905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_683 = _RAND_906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_684 = _RAND_907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_685 = _RAND_908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_686 = _RAND_909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_687 = _RAND_910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_688 = _RAND_911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_689 = _RAND_912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_690 = _RAND_913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_691 = _RAND_914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_692 = _RAND_915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_693 = _RAND_916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_694 = _RAND_917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_695 = _RAND_918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_696 = _RAND_919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_697 = _RAND_920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_698 = _RAND_921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_699 = _RAND_922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_700 = _RAND_923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_701 = _RAND_924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_702 = _RAND_925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_703 = _RAND_926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_704 = _RAND_927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_705 = _RAND_928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_706 = _RAND_929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_707 = _RAND_930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_708 = _RAND_931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_709 = _RAND_932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_710 = _RAND_933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_711 = _RAND_934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_712 = _RAND_935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_713 = _RAND_936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_714 = _RAND_937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_715 = _RAND_938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_716 = _RAND_939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_717 = _RAND_940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_718 = _RAND_941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_719 = _RAND_942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_720 = _RAND_943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_721 = _RAND_944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_722 = _RAND_945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_723 = _RAND_946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_724 = _RAND_947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_725 = _RAND_948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_726 = _RAND_949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_727 = _RAND_950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_728 = _RAND_951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_729 = _RAND_952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_730 = _RAND_953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_731 = _RAND_954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_732 = _RAND_955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_733 = _RAND_956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_734 = _RAND_957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_735 = _RAND_958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_736 = _RAND_959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_737 = _RAND_960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_738 = _RAND_961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_739 = _RAND_962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_740 = _RAND_963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_741 = _RAND_964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_742 = _RAND_965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_743 = _RAND_966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_744 = _RAND_967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_745 = _RAND_968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_746 = _RAND_969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_747 = _RAND_970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_748 = _RAND_971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_749 = _RAND_972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_750 = _RAND_973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_751 = _RAND_974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_752 = _RAND_975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_753 = _RAND_976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_754 = _RAND_977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_755 = _RAND_978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_756 = _RAND_979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_757 = _RAND_980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_758 = _RAND_981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_759 = _RAND_982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_760 = _RAND_983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_761 = _RAND_984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_762 = _RAND_985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_763 = _RAND_986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_764 = _RAND_987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_765 = _RAND_988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_766 = _RAND_989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_767 = _RAND_990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_768 = _RAND_991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_769 = _RAND_992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_770 = _RAND_993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_771 = _RAND_994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_772 = _RAND_995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_773 = _RAND_996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_774 = _RAND_997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_775 = _RAND_998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_776 = _RAND_999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_777 = _RAND_1000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_778 = _RAND_1001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_779 = _RAND_1002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_780 = _RAND_1003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_781 = _RAND_1004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_782 = _RAND_1005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_783 = _RAND_1006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_784 = _RAND_1007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_785 = _RAND_1008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_786 = _RAND_1009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_787 = _RAND_1010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_788 = _RAND_1011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_789 = _RAND_1012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_790 = _RAND_1013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_791 = _RAND_1014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_792 = _RAND_1015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_793 = _RAND_1016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_794 = _RAND_1017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_795 = _RAND_1018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_796 = _RAND_1019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_797 = _RAND_1020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_798 = _RAND_1021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_799 = _RAND_1022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_800 = _RAND_1023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_801 = _RAND_1024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 8'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    _T_132_re <= io_dIn_re;
    _T_132_im <= io_dIn_im;
    _T_133_re <= _T_132_re;
    _T_133_im <= _T_132_im;
    _T_134_re <= _T_133_re;
    _T_134_im <= _T_133_im;
    _T_135_re <= _T_134_re;
    _T_135_im <= _T_134_im;
    _T_136_re <= _T_135_re;
    _T_136_im <= _T_135_im;
    _T_137_re <= _T_136_re;
    _T_137_im <= _T_136_im;
    _T_138_re <= _T_137_re;
    _T_138_im <= _T_137_im;
    _T_139_re <= _T_138_re;
    _T_139_im <= _T_138_im;
    _T_140_re <= _T_139_re;
    _T_140_im <= _T_139_im;
    _T_141_re <= _T_140_re;
    _T_141_im <= _T_140_im;
    _T_142_re <= _T_141_re;
    _T_142_im <= _T_141_im;
    _T_143_re <= _T_142_re;
    _T_143_im <= _T_142_im;
    _T_144_re <= _T_143_re;
    _T_144_im <= _T_143_im;
    _T_145_re <= _T_144_re;
    _T_145_im <= _T_144_im;
    _T_146_re <= _T_145_re;
    _T_146_im <= _T_145_im;
    _T_147_re <= _T_146_re;
    _T_147_im <= _T_146_im;
    _T_148_re <= _T_147_re;
    _T_148_im <= _T_147_im;
    _T_149_re <= _T_148_re;
    _T_149_im <= _T_148_im;
    _T_150_re <= _T_149_re;
    _T_150_im <= _T_149_im;
    _T_151_re <= _T_150_re;
    _T_151_im <= _T_150_im;
    _T_152_re <= _T_151_re;
    _T_152_im <= _T_151_im;
    _T_153_re <= _T_152_re;
    _T_153_im <= _T_152_im;
    _T_154_re <= _T_153_re;
    _T_154_im <= _T_153_im;
    _T_155_re <= _T_154_re;
    _T_155_im <= _T_154_im;
    _T_156_re <= _T_155_re;
    _T_156_im <= _T_155_im;
    _T_157_re <= _T_156_re;
    _T_157_im <= _T_156_im;
    _T_158_re <= _T_157_re;
    _T_158_im <= _T_157_im;
    _T_159_re <= _T_158_re;
    _T_159_im <= _T_158_im;
    _T_160_re <= _T_159_re;
    _T_160_im <= _T_159_im;
    _T_161_re <= _T_160_re;
    _T_161_im <= _T_160_im;
    _T_162_re <= _T_161_re;
    _T_162_im <= _T_161_im;
    _T_163_re <= _T_162_re;
    _T_163_im <= _T_162_im;
    _T_164_re <= _T_163_re;
    _T_164_im <= _T_163_im;
    _T_165_re <= _T_164_re;
    _T_165_im <= _T_164_im;
    _T_166_re <= _T_165_re;
    _T_166_im <= _T_165_im;
    _T_167_re <= _T_166_re;
    _T_167_im <= _T_166_im;
    _T_168_re <= _T_167_re;
    _T_168_im <= _T_167_im;
    _T_169_re <= _T_168_re;
    _T_169_im <= _T_168_im;
    _T_170_re <= _T_169_re;
    _T_170_im <= _T_169_im;
    _T_171_re <= _T_170_re;
    _T_171_im <= _T_170_im;
    _T_172_re <= _T_171_re;
    _T_172_im <= _T_171_im;
    _T_173_re <= _T_172_re;
    _T_173_im <= _T_172_im;
    _T_174_re <= _T_173_re;
    _T_174_im <= _T_173_im;
    _T_175_re <= _T_174_re;
    _T_175_im <= _T_174_im;
    _T_176_re <= _T_175_re;
    _T_176_im <= _T_175_im;
    _T_177_re <= _T_176_re;
    _T_177_im <= _T_176_im;
    _T_178_re <= _T_177_re;
    _T_178_im <= _T_177_im;
    _T_179_re <= _T_178_re;
    _T_179_im <= _T_178_im;
    _T_180_re <= _T_179_re;
    _T_180_im <= _T_179_im;
    _T_181_re <= _T_180_re;
    _T_181_im <= _T_180_im;
    _T_182_re <= _T_181_re;
    _T_182_im <= _T_181_im;
    _T_183_re <= _T_182_re;
    _T_183_im <= _T_182_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_261_re <= Butterfly_io_out2_re;
    _T_261_im <= Butterfly_io_out2_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_329_re <= Switch_io_out1_re;
    _T_329_im <= Switch_io_out1_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_394_re <= Butterfly_1_io_out2_re;
    _T_394_im <= Butterfly_1_io_out2_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_402_re <= _T_401_re;
    _T_402_im <= _T_401_im;
    _T_403_re <= _T_402_re;
    _T_403_im <= _T_402_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_406_re <= _T_405_re;
    _T_406_im <= _T_405_im;
    _T_407_re <= _T_406_re;
    _T_407_im <= _T_406_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_409_re <= _T_408_re;
    _T_409_im <= _T_408_im;
    _T_410_re <= _T_409_re;
    _T_410_im <= _T_409_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_430_re <= Switch_1_io_out1_re;
    _T_430_im <= Switch_1_io_out1_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_463_re <= Butterfly_2_io_out2_re;
    _T_463_im <= Butterfly_2_io_out2_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_483_re <= Switch_2_io_out1_re;
    _T_483_im <= Switch_2_io_out1_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_500_re <= Butterfly_3_io_out2_re;
    _T_500_im <= Butterfly_3_io_out2_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_512_re <= Switch_3_io_out1_re;
    _T_512_im <= Switch_3_io_out1_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_521_re <= Butterfly_4_io_out2_re;
    _T_521_im <= Butterfly_4_io_out2_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_529_re <= Switch_4_io_out1_re;
    _T_529_im <= Switch_4_io_out1_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_534_re <= Butterfly_5_io_out2_re;
    _T_534_im <= Butterfly_5_io_out2_im;
    _T_535_re <= _T_534_re;
    _T_535_im <= _T_534_im;
    _T_540_re <= Switch_5_io_out1_re;
    _T_540_im <= Switch_5_io_out1_im;
    _T_541_re <= _T_540_re;
    _T_541_im <= _T_540_im;
    _T_543_re <= Butterfly_6_io_out2_re;
    _T_543_im <= Butterfly_6_io_out2_im;
    out1D1_re <= Switch_6_io_out1_re;
    out1D1_im <= Switch_6_io_out1_im;
    _T_544_re <= ComplexAdd_io_res_re;
    _T_544_im <= ComplexAdd_io_res_im;
    _T_545_re <= ComplexSub_io_res_re;
    _T_545_im <= ComplexSub_io_res_im;
    _T_546 <= io_din_valid;
    _T_547 <= _T_546;
    _T_548 <= _T_547;
    _T_549 <= _T_548;
    _T_550 <= _T_549;
    _T_551 <= _T_550;
    _T_552 <= _T_551;
    _T_553 <= _T_552;
    _T_554 <= _T_553;
    _T_555 <= _T_554;
    _T_556 <= _T_555;
    _T_557 <= _T_556;
    _T_558 <= _T_557;
    _T_559 <= _T_558;
    _T_560 <= _T_559;
    _T_561 <= _T_560;
    _T_562 <= _T_561;
    _T_563 <= _T_562;
    _T_564 <= _T_563;
    _T_565 <= _T_564;
    _T_566 <= _T_565;
    _T_567 <= _T_566;
    _T_568 <= _T_567;
    _T_569 <= _T_568;
    _T_570 <= _T_569;
    _T_571 <= _T_570;
    _T_572 <= _T_571;
    _T_573 <= _T_572;
    _T_574 <= _T_573;
    _T_575 <= _T_574;
    _T_576 <= _T_575;
    _T_577 <= _T_576;
    _T_578 <= _T_577;
    _T_579 <= _T_578;
    _T_580 <= _T_579;
    _T_581 <= _T_580;
    _T_582 <= _T_581;
    _T_583 <= _T_582;
    _T_584 <= _T_583;
    _T_585 <= _T_584;
    _T_586 <= _T_585;
    _T_587 <= _T_586;
    _T_588 <= _T_587;
    _T_589 <= _T_588;
    _T_590 <= _T_589;
    _T_591 <= _T_590;
    _T_592 <= _T_591;
    _T_593 <= _T_592;
    _T_594 <= _T_593;
    _T_595 <= _T_594;
    _T_596 <= _T_595;
    _T_597 <= _T_596;
    _T_598 <= _T_597;
    _T_599 <= _T_598;
    _T_600 <= _T_599;
    _T_601 <= _T_600;
    _T_602 <= _T_601;
    _T_603 <= _T_602;
    _T_604 <= _T_603;
    _T_605 <= _T_604;
    _T_606 <= _T_605;
    _T_607 <= _T_606;
    _T_608 <= _T_607;
    _T_609 <= _T_608;
    _T_610 <= _T_609;
    _T_611 <= _T_610;
    _T_612 <= _T_611;
    _T_613 <= _T_612;
    _T_614 <= _T_613;
    _T_615 <= _T_614;
    _T_616 <= _T_615;
    _T_617 <= _T_616;
    _T_618 <= _T_617;
    _T_619 <= _T_618;
    _T_620 <= _T_619;
    _T_621 <= _T_620;
    _T_622 <= _T_621;
    _T_623 <= _T_622;
    _T_624 <= _T_623;
    _T_625 <= _T_624;
    _T_626 <= _T_625;
    _T_627 <= _T_626;
    _T_628 <= _T_627;
    _T_629 <= _T_628;
    _T_630 <= _T_629;
    _T_631 <= _T_630;
    _T_632 <= _T_631;
    _T_633 <= _T_632;
    _T_634 <= _T_633;
    _T_635 <= _T_634;
    _T_636 <= _T_635;
    _T_637 <= _T_636;
    _T_638 <= _T_637;
    _T_639 <= _T_638;
    _T_640 <= _T_639;
    _T_641 <= _T_640;
    _T_642 <= _T_641;
    _T_643 <= _T_642;
    _T_644 <= _T_643;
    _T_645 <= _T_644;
    _T_646 <= _T_645;
    _T_647 <= _T_646;
    _T_648 <= _T_647;
    _T_649 <= _T_648;
    _T_650 <= _T_649;
    _T_651 <= _T_650;
    _T_652 <= _T_651;
    _T_653 <= _T_652;
    _T_654 <= _T_653;
    _T_655 <= _T_654;
    _T_656 <= _T_655;
    _T_657 <= _T_656;
    _T_658 <= _T_657;
    _T_659 <= _T_658;
    _T_660 <= _T_659;
    _T_661 <= _T_660;
    _T_662 <= _T_661;
    _T_663 <= _T_662;
    _T_664 <= _T_663;
    _T_665 <= _T_664;
    _T_666 <= _T_665;
    _T_667 <= _T_666;
    _T_668 <= _T_667;
    _T_669 <= _T_668;
    _T_670 <= _T_669;
    _T_671 <= _T_670;
    _T_672 <= _T_671;
    _T_673 <= _T_672;
    _T_674 <= _T_673;
    _T_675 <= _T_674;
    _T_676 <= _T_675;
    _T_677 <= _T_676;
    _T_678 <= _T_677;
    _T_679 <= _T_678;
    _T_680 <= _T_679;
    _T_681 <= _T_680;
    _T_682 <= _T_681;
    _T_683 <= _T_682;
    _T_684 <= _T_683;
    _T_685 <= _T_684;
    _T_686 <= _T_685;
    _T_687 <= _T_686;
    _T_688 <= _T_687;
    _T_689 <= _T_688;
    _T_690 <= _T_689;
    _T_691 <= _T_690;
    _T_692 <= _T_691;
    _T_693 <= _T_692;
    _T_694 <= _T_693;
    _T_695 <= _T_694;
    _T_696 <= _T_695;
    _T_697 <= _T_696;
    _T_698 <= _T_697;
    _T_699 <= _T_698;
    _T_700 <= _T_699;
    _T_701 <= _T_700;
    _T_702 <= _T_701;
    _T_703 <= _T_702;
    _T_704 <= _T_703;
    _T_705 <= _T_704;
    _T_706 <= _T_705;
    _T_707 <= _T_706;
    _T_708 <= _T_707;
    _T_709 <= _T_708;
    _T_710 <= _T_709;
    _T_711 <= _T_710;
    _T_712 <= _T_711;
    _T_713 <= _T_712;
    _T_714 <= _T_713;
    _T_715 <= _T_714;
    _T_716 <= _T_715;
    _T_717 <= _T_716;
    _T_718 <= _T_717;
    _T_719 <= _T_718;
    _T_720 <= _T_719;
    _T_721 <= _T_720;
    _T_722 <= _T_721;
    _T_723 <= _T_722;
    _T_724 <= _T_723;
    _T_725 <= _T_724;
    _T_726 <= _T_725;
    _T_727 <= _T_726;
    _T_728 <= _T_727;
    _T_729 <= _T_728;
    _T_730 <= _T_729;
    _T_731 <= _T_730;
    _T_732 <= _T_731;
    _T_733 <= _T_732;
    _T_734 <= _T_733;
    _T_735 <= _T_734;
    _T_736 <= _T_735;
    _T_737 <= _T_736;
    _T_738 <= _T_737;
    _T_739 <= _T_738;
    _T_740 <= _T_739;
    _T_741 <= _T_740;
    _T_742 <= _T_741;
    _T_743 <= _T_742;
    _T_744 <= _T_743;
    _T_745 <= _T_744;
    _T_746 <= _T_745;
    _T_747 <= _T_746;
    _T_748 <= _T_747;
    _T_749 <= _T_748;
    _T_750 <= _T_749;
    _T_751 <= _T_750;
    _T_752 <= _T_751;
    _T_753 <= _T_752;
    _T_754 <= _T_753;
    _T_755 <= _T_754;
    _T_756 <= _T_755;
    _T_757 <= _T_756;
    _T_758 <= _T_757;
    _T_759 <= _T_758;
    _T_760 <= _T_759;
    _T_761 <= _T_760;
    _T_762 <= _T_761;
    _T_763 <= _T_762;
    _T_764 <= _T_763;
    _T_765 <= _T_764;
    _T_766 <= _T_765;
    _T_767 <= _T_766;
    _T_768 <= _T_767;
    _T_769 <= _T_768;
    _T_770 <= _T_769;
    _T_771 <= _T_770;
    _T_772 <= _T_771;
    _T_773 <= _T_772;
    _T_774 <= _T_773;
    _T_775 <= _T_774;
    _T_776 <= _T_775;
    _T_777 <= _T_776;
    _T_778 <= _T_777;
    _T_779 <= _T_778;
    _T_780 <= _T_779;
    _T_781 <= _T_780;
    _T_782 <= _T_781;
    _T_783 <= _T_782;
    _T_784 <= _T_783;
    _T_785 <= _T_784;
    _T_786 <= _T_785;
    _T_787 <= _T_786;
    _T_788 <= _T_787;
    _T_789 <= _T_788;
    _T_790 <= _T_789;
    _T_791 <= _T_790;
    _T_792 <= _T_791;
    _T_793 <= _T_792;
    _T_794 <= _T_793;
    _T_795 <= _T_794;
    _T_796 <= _T_795;
    _T_797 <= _T_796;
    _T_798 <= _T_797;
    _T_799 <= _T_798;
    _T_800 <= _T_799;
    _T_801 <= _T_800;
  end
endmodule
