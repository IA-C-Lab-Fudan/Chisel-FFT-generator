module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T; // @[Butterfly.scala 57:28]
  wire [63:0] _T_1; // @[Butterfly.scala 57:52]
  wire [63:0] _T_4; // @[Butterfly.scala 57:40]
  wire [63:0] _T_5; // @[Butterfly.scala 58:28]
  wire [63:0] _T_6; // @[Butterfly.scala 58:52]
  wire [63:0] _T_9; // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2; // @[Butterfly.scala 58:15]
  assign _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  assign _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  assign _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  assign _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  assign _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  assign _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  assign _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT2048RAM(
    input clk_in1_p,
    input clk_in1_n,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
    wire clock;
    clk_wiz_0 clk_wiz_0_inst0
       (
        // Clock out ports
        .clk_out1(clock),     // output clk_out1
       // Clock in ports
        .clk_in1_p(clk_in1_p),    // input clk_in1_p
        .clk_in1_n(clk_in1_n));    // input clk_in1_n
  wire  BRAM_clock; // @[FFT.scala 62:23]
  wire  BRAM_en; // @[FFT.scala 62:23]
  wire [9:0] BRAM_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_1_clock; // @[FFT.scala 62:23]
  wire  BRAM_1_en; // @[FFT.scala 62:23]
  wire [8:0] BRAM_1_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_1_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_2_clock; // @[FFT.scala 62:23]
  wire  BRAM_2_en; // @[FFT.scala 62:23]
  wire [7:0] BRAM_2_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_2_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_3_clock; // @[FFT.scala 62:23]
  wire  BRAM_3_en; // @[FFT.scala 62:23]
  wire [6:0] BRAM_3_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_3_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_4_clock; // @[FFT.scala 62:23]
  wire  BRAM_4_en; // @[FFT.scala 62:23]
  wire [5:0] BRAM_4_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_4_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_5_clock; // @[FFT.scala 62:23]
  wire  BRAM_5_en; // @[FFT.scala 62:23]
  wire [4:0] BRAM_5_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_5_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_8_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_8_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_8_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_8_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_8_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_9_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_9_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_9_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_9_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_9_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [10:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [10:0] _T_1; // @[FFT.scala 42:16]
  reg [10:0] cntD1; // @[FFT.scala 44:22]
  reg [31:0] _RAND_1;
  reg [10:0] cntD2; // @[FFT.scala 45:22]
  reg [31:0] _RAND_2;
  reg [31:0] out1_0_re; // @[FFT.scala 50:23]
  reg [31:0] _RAND_3;
  reg [31:0] out1_0_im; // @[FFT.scala 50:23]
  reg [31:0] _RAND_4;
  reg [31:0] out2_0_re; // @[FFT.scala 51:23]
  reg [31:0] _RAND_5;
  reg [31:0] out2_0_im; // @[FFT.scala 51:23]
  reg [31:0] _RAND_6;
  wire [63:0] _T_176;
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [31:0] _T_393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [31:0] _T_402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [31:0] _T_406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [31:0] _T_409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [31:0] _T_409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_521;
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_522;
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_523;
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_524;
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_525;
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_526;
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_527;
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_528;
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_529;
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_530;
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_531;
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_532;
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_533;
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_534;
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_535;
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_536;
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_537;
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_538;
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_539;
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_540;
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_541;
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_552;
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_553;
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_554;
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_557;
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_558;
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_559;
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_560;
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_561;
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_562;
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_563;
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_564;
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_565;
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_566;
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_567;
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_568;
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_569;
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_570;
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_571;
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_572;
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_573;
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_574;
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_575;
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_576;
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_577;
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_578;
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_579;
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_580;
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_581;
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_582;
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_583;
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_584;
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_585;
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_586;
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_587;
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_588;
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_589;
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_590;
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_591;
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_592;
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_593;
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_594;
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_595;
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_596;
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_597;
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_598;
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_599;
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_600;
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_601;
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_602;
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_603;
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_604;
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_605;
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_606;
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_607;
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_608;
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_609;
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_610;
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_611;
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_612;
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_613;
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_614;
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_615;
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_616;
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_617;
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_618;
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_619;
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_620;
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_621;
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_622;
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_623;
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_624;
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_625;
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_626;
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_627;
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_628;
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_629;
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_630;
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_631;
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_632;
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_633;
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_634;
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_635;
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_636;
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_637;
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_638;
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_639;
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_640;
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_641;
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_642;
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_643;
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_644;
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_645;
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_646;
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_647;
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_648;
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_649;
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_650;
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_651;
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_652;
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_653;
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_654;
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_655;
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_656;
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_657;
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_658;
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_659;
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_660;
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_661;
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_662;
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_663;
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_664;
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_665;
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_666;
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_667;
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_668;
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_669;
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_670;
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_671;
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_672;
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_673;
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_674;
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_675;
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_676;
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_677;
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_678;
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_679;
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_680;
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_681;
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_682;
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_683;
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_684;
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_685;
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_686;
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_687;
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_688;
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_689;
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_690;
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_691;
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_692;
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_693;
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_694;
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_695;
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_696;
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_697;
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_698;
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_699;
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_700;
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_701;
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_702;
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_703;
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_704;
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_705;
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_706;
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_707;
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_708;
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_709;
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_710;
  reg [31:0] _T_533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_711;
  reg [31:0] _T_533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_712;
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_713;
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_714;
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_715;
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_716;
  reg [31:0] _T_536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_717;
  reg [31:0] _T_536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_718;
  reg [31:0] _T_537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_719;
  reg [31:0] _T_537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_720;
  reg [31:0] _T_538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_721;
  reg [31:0] _T_538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_722;
  reg [31:0] _T_539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_723;
  reg [31:0] _T_539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_724;
  reg [31:0] _T_540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_725;
  reg [31:0] _T_540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_726;
  reg [31:0] _T_541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_727;
  reg [31:0] _T_541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_728;
  reg [31:0] _T_542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_729;
  reg [31:0] _T_542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_730;
  reg [31:0] _T_543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_731;
  reg [31:0] _T_543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_732;
  reg [31:0] _T_544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_733;
  reg [31:0] _T_544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_734;
  reg [31:0] _T_545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_735;
  reg [31:0] _T_545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_736;
  reg [31:0] _T_546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_737;
  reg [31:0] _T_546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_738;
  reg [31:0] _T_547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_739;
  reg [31:0] _T_547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_740;
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_741;
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_742;
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_743;
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_744;
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_745;
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_746;
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_747;
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_748;
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_749;
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_750;
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_751;
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_752;
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_753;
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_754;
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_755;
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_756;
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_757;
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_758;
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_759;
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_760;
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_761;
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_762;
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_763;
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_764;
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_765;
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_766;
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_767;
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_768;
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_769;
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_771;
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_772;
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_773;
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_781;
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_782;
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_783;
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_784;
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_785;
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_786;
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_787;
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_788;
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_789;
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_790;
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_791;
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_792;
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_793;
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_794;
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_795;
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_796;
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_797;
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_798;
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_799;
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_800;
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_801;
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_802;
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_803;
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_804;
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_805;
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_806;
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_807;
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_808;
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_809;
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_810;
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_811;
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_812;
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_813;
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_814;
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_815;
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_816;
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_817;
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_818;
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_819;
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_820;
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_821;
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_822;
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_823;
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_824;
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_825;
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_826;
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_827;
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_828;
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_829;
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_830;
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_831;
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_832;
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_833;
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_834;
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_835;
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_836;
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_837;
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_838;
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_839;
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_840;
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_841;
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_842;
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_843;
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_844;
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_845;
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_846;
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_847;
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_848;
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_849;
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_850;
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_851;
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_852;
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_853;
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_854;
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_855;
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_856;
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_857;
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_858;
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_859;
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_860;
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_861;
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_862;
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_863;
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_864;
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_865;
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_866;
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_867;
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_868;
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_869;
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_870;
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_871;
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_872;
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_873;
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_874;
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_875;
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_876;
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_877;
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_878;
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_879;
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_880;
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_881;
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_882;
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_883;
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_884;
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_885;
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_886;
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_887;
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_888;
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_889;
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_890;
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_891;
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_892;
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_893;
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_894;
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_895;
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_896;
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_897;
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_898;
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_899;
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_900;
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_901;
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_902;
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_903;
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_904;
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_905;
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_906;
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_907;
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_908;
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_909;
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_910;
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_911;
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_912;
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_913;
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_914;
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_915;
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_916;
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_917;
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_918;
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_919;
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_920;
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_921;
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_922;
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_923;
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_924;
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_925;
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_926;
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_927;
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_928;
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_929;
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_930;
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_931;
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_932;
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_933;
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_934;
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_935;
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_936;
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_937;
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_938;
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_939;
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_940;
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_941;
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_942;
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_943;
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_944;
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_945;
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_946;
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_947;
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_948;
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_949;
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_950;
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_951;
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_952;
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_953;
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_954;
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_955;
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_956;
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_957;
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_958;
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_959;
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_960;
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_961;
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_962;
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_963;
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_964;
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_965;
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_966;
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_967;
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_968;
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_969;
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_970;
  reg [31:0] _T_663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_971;
  reg [31:0] _T_663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_972;
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_973;
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_974;
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_975;
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_976;
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_977;
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_978;
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_979;
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_980;
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_981;
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_982;
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_983;
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_984;
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_985;
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_986;
  reg [31:0] _T_671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_987;
  reg [31:0] _T_671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_988;
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_989;
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_990;
  reg [31:0] _T_673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_991;
  reg [31:0] _T_673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_992;
  reg [31:0] _T_674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_993;
  reg [31:0] _T_674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_994;
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_995;
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_996;
  reg [31:0] _T_676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_997;
  reg [31:0] _T_676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_998;
  reg [31:0] _T_677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_999;
  reg [31:0] _T_677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1000;
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1001;
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1002;
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1003;
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1004;
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1005;
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1006;
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1007;
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1008;
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1009;
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1010;
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1011;
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1012;
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1013;
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1014;
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1015;
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1016;
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1017;
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1018;
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1019;
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1020;
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1021;
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1022;
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1023;
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1024;
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1025;
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1026;
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1027;
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1028;
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1029;
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1030;
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1031;
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1032;
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1033;
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1034;
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1035;
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1036;
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1037;
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1038;
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1039;
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1040;
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1041;
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1042;
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1043;
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1044;
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1045;
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1046;
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1047;
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1048;
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1049;
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1050;
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1051;
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1052;
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1053;
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1054;
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1055;
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1056;
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1057;
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1058;
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1059;
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1060;
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1061;
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1062;
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1063;
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1064;
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1065;
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1066;
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1067;
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1068;
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1069;
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1070;
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1071;
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1072;
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1073;
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1074;
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1075;
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1076;
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1077;
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1078;
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1079;
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1080;
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1081;
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1082;
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1083;
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1084;
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1085;
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1086;
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1087;
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1088;
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1089;
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1090;
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1091;
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1092;
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1093;
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1094;
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1095;
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1096;
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1097;
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1098;
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1099;
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1100;
  reg [31:0] _T_728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1101;
  reg [31:0] _T_728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1102;
  reg [31:0] _T_729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1103;
  reg [31:0] _T_729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1104;
  reg [31:0] _T_730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1105;
  reg [31:0] _T_730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1106;
  reg [31:0] _T_731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1107;
  reg [31:0] _T_731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1108;
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1109;
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1110;
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1111;
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1112;
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1113;
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1114;
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1115;
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1116;
  reg [31:0] _T_736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1117;
  reg [31:0] _T_736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1118;
  reg [31:0] _T_737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1119;
  reg [31:0] _T_737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1120;
  reg [31:0] _T_738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1121;
  reg [31:0] _T_738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1122;
  reg [31:0] _T_739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1123;
  reg [31:0] _T_739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1124;
  reg [31:0] _T_740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1125;
  reg [31:0] _T_740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1126;
  reg [31:0] _T_741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1127;
  reg [31:0] _T_741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1128;
  reg [31:0] _T_742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1129;
  reg [31:0] _T_742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1130;
  reg [31:0] _T_743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1131;
  reg [31:0] _T_743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1132;
  reg [31:0] _T_744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1133;
  reg [31:0] _T_744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1134;
  reg [31:0] _T_745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1135;
  reg [31:0] _T_745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1136;
  reg [31:0] _T_746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1137;
  reg [31:0] _T_746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1138;
  reg [31:0] _T_747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1139;
  reg [31:0] _T_747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1140;
  reg [31:0] _T_748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1141;
  reg [31:0] _T_748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1142;
  reg [31:0] _T_749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1143;
  reg [31:0] _T_749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1144;
  reg [31:0] _T_750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1145;
  reg [31:0] _T_750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1146;
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1147;
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1148;
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1149;
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1150;
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1151;
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1152;
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1153;
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1154;
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1155;
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1156;
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1157;
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1158;
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1159;
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1160;
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1161;
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1162;
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1163;
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1164;
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1165;
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1166;
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1167;
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1168;
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1169;
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1170;
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1171;
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1172;
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1173;
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1174;
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1175;
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1176;
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1177;
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1178;
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1179;
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1180;
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1181;
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1182;
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1183;
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1184;
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1185;
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1186;
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1187;
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1188;
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1189;
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1190;
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1191;
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1192;
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1193;
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1194;
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1195;
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1196;
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1197;
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1198;
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1199;
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1200;
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1201;
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1202;
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1203;
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1204;
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1205;
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1206;
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1207;
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1208;
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1209;
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1210;
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1211;
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1212;
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1213;
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1214;
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1215;
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1216;
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1217;
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1218;
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1219;
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1220;
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1221;
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1222;
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1223;
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1224;
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1225;
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1226;
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1227;
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1228;
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1229;
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1230;
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1231;
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1232;
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1233;
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1234;
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1235;
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1236;
  reg [31:0] _T_796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1237;
  reg [31:0] _T_796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1238;
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1239;
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1240;
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1241;
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1242;
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1243;
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1244;
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1245;
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1246;
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1247;
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1248;
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1249;
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1250;
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1251;
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1252;
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1253;
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1254;
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1255;
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1256;
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1257;
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1258;
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1259;
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1260;
  reg [31:0] _T_808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1261;
  reg [31:0] _T_808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1262;
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1263;
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1264;
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1265;
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1266;
  reg [31:0] _T_811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1267;
  reg [31:0] _T_811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1268;
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1269;
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1270;
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1271;
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1272;
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1273;
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1274;
  reg [31:0] _T_815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1275;
  reg [31:0] _T_815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1276;
  reg [31:0] _T_816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1277;
  reg [31:0] _T_816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1278;
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1279;
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1280;
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1281;
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1282;
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1283;
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1284;
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1285;
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1286;
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1287;
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1288;
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1289;
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1290;
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1291;
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1292;
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1293;
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1294;
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1295;
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1296;
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1297;
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1298;
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1299;
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1300;
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1301;
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1302;
  reg [31:0] _T_829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1303;
  reg [31:0] _T_829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1304;
  reg [31:0] _T_830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1305;
  reg [31:0] _T_830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1306;
  reg [31:0] _T_831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1307;
  reg [31:0] _T_831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1308;
  reg [31:0] _T_832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1309;
  reg [31:0] _T_832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1310;
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1311;
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1312;
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1313;
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1314;
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1315;
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1316;
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1317;
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1318;
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1319;
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1320;
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1321;
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1322;
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1323;
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1324;
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1325;
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1326;
  reg [31:0] _T_841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1327;
  reg [31:0] _T_841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1328;
  reg [31:0] _T_842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1329;
  reg [31:0] _T_842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1330;
  reg [31:0] _T_843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1331;
  reg [31:0] _T_843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1332;
  reg [31:0] _T_844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1333;
  reg [31:0] _T_844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1334;
  reg [31:0] _T_845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1335;
  reg [31:0] _T_845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1336;
  reg [31:0] _T_846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1337;
  reg [31:0] _T_846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1338;
  reg [31:0] _T_847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1339;
  reg [31:0] _T_847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1340;
  reg [31:0] _T_848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1341;
  reg [31:0] _T_848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1342;
  reg [31:0] _T_849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1343;
  reg [31:0] _T_849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1344;
  reg [31:0] _T_850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1345;
  reg [31:0] _T_850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1346;
  reg [31:0] _T_851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1347;
  reg [31:0] _T_851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1348;
  reg [31:0] _T_852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1349;
  reg [31:0] _T_852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1350;
  reg [31:0] _T_853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1351;
  reg [31:0] _T_853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1352;
  reg [31:0] _T_854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1353;
  reg [31:0] _T_854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1354;
  reg [31:0] _T_855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1355;
  reg [31:0] _T_855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1356;
  reg [31:0] _T_856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1357;
  reg [31:0] _T_856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1358;
  reg [31:0] _T_857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1359;
  reg [31:0] _T_857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1360;
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1361;
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1362;
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1363;
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1364;
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1365;
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1366;
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1367;
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1368;
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1369;
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1370;
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1371;
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1372;
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1373;
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1374;
  reg [31:0] _T_865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1375;
  reg [31:0] _T_865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1376;
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1377;
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1378;
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1379;
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1380;
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1381;
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1382;
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1383;
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1384;
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1385;
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1386;
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1387;
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1388;
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1389;
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1390;
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1391;
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1392;
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1393;
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1394;
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1395;
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1396;
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1397;
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1398;
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1399;
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1400;
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1401;
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1402;
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1403;
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1404;
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1405;
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1406;
  reg [31:0] _T_881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1407;
  reg [31:0] _T_881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1408;
  reg [31:0] _T_882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1409;
  reg [31:0] _T_882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1410;
  reg [31:0] _T_883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1411;
  reg [31:0] _T_883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1412;
  reg [31:0] _T_884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1413;
  reg [31:0] _T_884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1414;
  reg [31:0] _T_885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1415;
  reg [31:0] _T_885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1416;
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1417;
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1418;
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1419;
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1420;
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1421;
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1422;
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1423;
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1424;
  reg [31:0] _T_890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1425;
  reg [31:0] _T_890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1426;
  reg [31:0] _T_891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1427;
  reg [31:0] _T_891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1428;
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1429;
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1430;
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1431;
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1432;
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1433;
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1434;
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1435;
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1436;
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1437;
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1438;
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1439;
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1440;
  reg [31:0] _T_898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1441;
  reg [31:0] _T_898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1442;
  reg [31:0] _T_899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1443;
  reg [31:0] _T_899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1444;
  reg [31:0] _T_900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1445;
  reg [31:0] _T_900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1446;
  reg [31:0] _T_901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1447;
  reg [31:0] _T_901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1448;
  reg [31:0] _T_902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1449;
  reg [31:0] _T_902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1450;
  reg [31:0] _T_903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1451;
  reg [31:0] _T_903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1452;
  reg [31:0] _T_904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1453;
  reg [31:0] _T_904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1454;
  reg [31:0] _T_905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1455;
  reg [31:0] _T_905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1456;
  reg [31:0] _T_906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1457;
  reg [31:0] _T_906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1458;
  reg [31:0] _T_907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1459;
  reg [31:0] _T_907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1460;
  reg [31:0] _T_908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1461;
  reg [31:0] _T_908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1462;
  reg [31:0] _T_909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1463;
  reg [31:0] _T_909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1464;
  reg [31:0] _T_910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1465;
  reg [31:0] _T_910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1466;
  reg [31:0] _T_911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1467;
  reg [31:0] _T_911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1468;
  reg [31:0] _T_912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1469;
  reg [31:0] _T_912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1470;
  reg [31:0] _T_913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1471;
  reg [31:0] _T_913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1472;
  reg [31:0] _T_914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1473;
  reg [31:0] _T_914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1474;
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1475;
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1476;
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1477;
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1478;
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1479;
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1480;
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1481;
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1482;
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1483;
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1484;
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1485;
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1486;
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1487;
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1488;
  reg [31:0] _T_922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1489;
  reg [31:0] _T_922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1490;
  reg [31:0] _T_923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1491;
  reg [31:0] _T_923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1492;
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1493;
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1494;
  reg [31:0] _T_925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1495;
  reg [31:0] _T_925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1496;
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1497;
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1498;
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1499;
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1500;
  reg [31:0] _T_928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1501;
  reg [31:0] _T_928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1502;
  reg [31:0] _T_929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1503;
  reg [31:0] _T_929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1504;
  reg [31:0] _T_930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1505;
  reg [31:0] _T_930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1506;
  reg [31:0] _T_931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1507;
  reg [31:0] _T_931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1508;
  reg [31:0] _T_932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1509;
  reg [31:0] _T_932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1510;
  reg [31:0] _T_933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1511;
  reg [31:0] _T_933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1512;
  reg [31:0] _T_934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1513;
  reg [31:0] _T_934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1514;
  reg [31:0] _T_935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1515;
  reg [31:0] _T_935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1516;
  reg [31:0] _T_936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1517;
  reg [31:0] _T_936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1518;
  reg [31:0] _T_937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1519;
  reg [31:0] _T_937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1520;
  reg [31:0] _T_938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1521;
  reg [31:0] _T_938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1522;
  reg [31:0] _T_939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1523;
  reg [31:0] _T_939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1524;
  reg [31:0] _T_940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1525;
  reg [31:0] _T_940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1526;
  reg [31:0] _T_941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1527;
  reg [31:0] _T_941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1528;
  reg [31:0] _T_942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1529;
  reg [31:0] _T_942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1530;
  reg [31:0] _T_943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1531;
  reg [31:0] _T_943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1532;
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1533;
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1534;
  reg [31:0] _T_945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1535;
  reg [31:0] _T_945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1536;
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1537;
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1538;
  reg [31:0] _T_947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1539;
  reg [31:0] _T_947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1540;
  reg [31:0] _T_948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1541;
  reg [31:0] _T_948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1542;
  reg [31:0] _T_949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1543;
  reg [31:0] _T_949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1544;
  reg [31:0] _T_950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1545;
  reg [31:0] _T_950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1546;
  reg [31:0] _T_951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1547;
  reg [31:0] _T_951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1548;
  reg [31:0] _T_952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1549;
  reg [31:0] _T_952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1550;
  reg [31:0] _T_953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1551;
  reg [31:0] _T_953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1552;
  reg [31:0] _T_954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1553;
  reg [31:0] _T_954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1554;
  reg [31:0] _T_955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1555;
  reg [31:0] _T_955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1556;
  reg [31:0] _T_956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1557;
  reg [31:0] _T_956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1558;
  reg [31:0] _T_957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1559;
  reg [31:0] _T_957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1560;
  reg [31:0] _T_958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1561;
  reg [31:0] _T_958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1562;
  reg [31:0] _T_959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1563;
  reg [31:0] _T_959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1564;
  reg [31:0] _T_960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1565;
  reg [31:0] _T_960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1566;
  reg [31:0] _T_961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1567;
  reg [31:0] _T_961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1568;
  reg [31:0] _T_962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1569;
  reg [31:0] _T_962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1570;
  reg [31:0] _T_963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1571;
  reg [31:0] _T_963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1572;
  reg [31:0] _T_964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1573;
  reg [31:0] _T_964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1574;
  reg [31:0] _T_965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1575;
  reg [31:0] _T_965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1576;
  reg [31:0] _T_966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1577;
  reg [31:0] _T_966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1578;
  reg [31:0] _T_967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1579;
  reg [31:0] _T_967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1580;
  reg [31:0] _T_968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1581;
  reg [31:0] _T_968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1582;
  reg [31:0] _T_969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1583;
  reg [31:0] _T_969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1584;
  reg [31:0] _T_970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1585;
  reg [31:0] _T_970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1586;
  reg [31:0] _T_971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1587;
  reg [31:0] _T_971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1588;
  reg [31:0] _T_972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1589;
  reg [31:0] _T_972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1590;
  reg [31:0] _T_973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1591;
  reg [31:0] _T_973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1592;
  reg [31:0] _T_974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1593;
  reg [31:0] _T_974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1594;
  reg [31:0] _T_975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1595;
  reg [31:0] _T_975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1596;
  reg [31:0] _T_976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1597;
  reg [31:0] _T_976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1598;
  reg [31:0] _T_977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1599;
  reg [31:0] _T_977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1600;
  reg [31:0] _T_978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1601;
  reg [31:0] _T_978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1602;
  reg [31:0] _T_979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1603;
  reg [31:0] _T_979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1604;
  reg [31:0] _T_980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1605;
  reg [31:0] _T_980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1606;
  reg [31:0] _T_981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1607;
  reg [31:0] _T_981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1608;
  reg [31:0] _T_982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1609;
  reg [31:0] _T_982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1610;
  reg [31:0] _T_983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1611;
  reg [31:0] _T_983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1612;
  reg [31:0] _T_984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1613;
  reg [31:0] _T_984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1614;
  reg [31:0] _T_985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1615;
  reg [31:0] _T_985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1616;
  reg [31:0] _T_986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1617;
  reg [31:0] _T_986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1618;
  reg [31:0] _T_987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1619;
  reg [31:0] _T_987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1620;
  reg [31:0] _T_988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1621;
  reg [31:0] _T_988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1622;
  reg [31:0] _T_989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1623;
  reg [31:0] _T_989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1624;
  reg [31:0] _T_990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1625;
  reg [31:0] _T_990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1626;
  reg [31:0] _T_991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1627;
  reg [31:0] _T_991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1628;
  reg [31:0] _T_992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1629;
  reg [31:0] _T_992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1630;
  reg [31:0] _T_993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1631;
  reg [31:0] _T_993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1632;
  reg [31:0] _T_994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1633;
  reg [31:0] _T_994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1634;
  reg [31:0] _T_995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1635;
  reg [31:0] _T_995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1636;
  reg [31:0] _T_996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1637;
  reg [31:0] _T_996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1638;
  reg [31:0] _T_997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1639;
  reg [31:0] _T_997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1640;
  reg [31:0] _T_998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1641;
  reg [31:0] _T_998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1642;
  reg [31:0] _T_999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1643;
  reg [31:0] _T_999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1644;
  reg [31:0] _T_1000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1645;
  reg [31:0] _T_1000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1646;
  reg [31:0] _T_1001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1647;
  reg [31:0] _T_1001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1648;
  reg [31:0] _T_1002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1649;
  reg [31:0] _T_1002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1650;
  reg [31:0] _T_1003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1651;
  reg [31:0] _T_1003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1652;
  reg [31:0] _T_1004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1653;
  reg [31:0] _T_1004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1654;
  reg [31:0] _T_1005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1655;
  reg [31:0] _T_1005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1656;
  reg [31:0] _T_1006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1657;
  reg [31:0] _T_1006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1658;
  reg [31:0] _T_1007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1659;
  reg [31:0] _T_1007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1660;
  reg [31:0] _T_1008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1661;
  reg [31:0] _T_1008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1662;
  reg [31:0] _T_1009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1663;
  reg [31:0] _T_1009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1664;
  reg [31:0] _T_1010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1665;
  reg [31:0] _T_1010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1666;
  reg [31:0] _T_1011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1667;
  reg [31:0] _T_1011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1668;
  reg [31:0] _T_1012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1669;
  reg [31:0] _T_1012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1670;
  reg [31:0] _T_1013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1671;
  reg [31:0] _T_1013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1672;
  reg [31:0] _T_1014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1673;
  reg [31:0] _T_1014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1674;
  reg [31:0] _T_1015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1675;
  reg [31:0] _T_1015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1676;
  reg [31:0] _T_1016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1677;
  reg [31:0] _T_1016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1678;
  reg [31:0] _T_1017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1679;
  reg [31:0] _T_1017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1680;
  reg [31:0] _T_1018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1681;
  reg [31:0] _T_1018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1682;
  reg [31:0] _T_1019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1683;
  reg [31:0] _T_1019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1684;
  reg [31:0] _T_1020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1685;
  reg [31:0] _T_1020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1686;
  reg [31:0] _T_1021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1687;
  reg [31:0] _T_1021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1688;
  reg [31:0] _T_1022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1689;
  reg [31:0] _T_1022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1690;
  reg [31:0] _T_1023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1691;
  reg [31:0] _T_1023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1692;
  reg [31:0] _T_1024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1693;
  reg [31:0] _T_1024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1694;
  reg [31:0] _T_1025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1695;
  reg [31:0] _T_1025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1696;
  reg [31:0] _T_1026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1697;
  reg [31:0] _T_1026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1698;
  reg [31:0] _T_1027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1699;
  reg [31:0] _T_1027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1700;
  reg [31:0] _T_1028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1701;
  reg [31:0] _T_1028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1702;
  reg [31:0] _T_1029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1703;
  reg [31:0] _T_1029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1704;
  reg [31:0] _T_1030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1705;
  reg [31:0] _T_1030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1706;
  reg [31:0] _T_1031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1707;
  reg [31:0] _T_1031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1708;
  reg [31:0] _T_1032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1709;
  reg [31:0] _T_1032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1710;
  reg [31:0] _T_1033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1711;
  reg [31:0] _T_1033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1712;
  reg [31:0] _T_1034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1713;
  reg [31:0] _T_1034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1714;
  reg [31:0] _T_1035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1715;
  reg [31:0] _T_1035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1716;
  reg [31:0] _T_1036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1717;
  reg [31:0] _T_1036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1718;
  reg [31:0] _T_1037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1719;
  reg [31:0] _T_1037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1720;
  reg [31:0] _T_1038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1721;
  reg [31:0] _T_1038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1722;
  reg [31:0] _T_1039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1723;
  reg [31:0] _T_1039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1724;
  reg [31:0] _T_1040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1725;
  reg [31:0] _T_1040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1726;
  reg [31:0] _T_1041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1727;
  reg [31:0] _T_1041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1728;
  reg [31:0] _T_1042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1729;
  reg [31:0] _T_1042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1730;
  reg [31:0] _T_1043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1731;
  reg [31:0] _T_1043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1732;
  reg [31:0] _T_1044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1733;
  reg [31:0] _T_1044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1734;
  reg [31:0] _T_1045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1735;
  reg [31:0] _T_1045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1736;
  reg [31:0] _T_1046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1737;
  reg [31:0] _T_1046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1738;
  reg [31:0] _T_1047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1739;
  reg [31:0] _T_1047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1740;
  reg [31:0] _T_1048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1741;
  reg [31:0] _T_1048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1742;
  reg [31:0] _T_1049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1743;
  reg [31:0] _T_1049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1744;
  reg [31:0] _T_1050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1745;
  reg [31:0] _T_1050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1746;
  reg [31:0] _T_1051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1747;
  reg [31:0] _T_1051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1748;
  reg [31:0] _T_1052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1749;
  reg [31:0] _T_1052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1750;
  reg [31:0] _T_1053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1751;
  reg [31:0] _T_1053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1752;
  reg [31:0] _T_1054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1753;
  reg [31:0] _T_1054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1754;
  reg [31:0] _T_1055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1755;
  reg [31:0] _T_1055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1756;
  reg [31:0] _T_1056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1757;
  reg [31:0] _T_1056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1758;
  reg [31:0] _T_1057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1759;
  reg [31:0] _T_1057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1760;
  reg [31:0] _T_1058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1761;
  reg [31:0] _T_1058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1762;
  reg [31:0] _T_1059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1763;
  reg [31:0] _T_1059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1764;
  reg [31:0] _T_1060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1765;
  reg [31:0] _T_1060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1766;
  reg [31:0] _T_1061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1767;
  reg [31:0] _T_1061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1768;
  reg [31:0] _T_1062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1769;
  reg [31:0] _T_1062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1770;
  reg [31:0] _T_1063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1771;
  reg [31:0] _T_1063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1772;
  reg [31:0] _T_1064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1773;
  reg [31:0] _T_1064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1774;
  reg [31:0] _T_1065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1775;
  reg [31:0] _T_1065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1776;
  reg [31:0] _T_1066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1777;
  reg [31:0] _T_1066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1778;
  reg [31:0] _T_1067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1779;
  reg [31:0] _T_1067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1780;
  reg [31:0] _T_1068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1781;
  reg [31:0] _T_1068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1782;
  reg [31:0] _T_1069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1783;
  reg [31:0] _T_1069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1784;
  reg [31:0] _T_1070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1785;
  reg [31:0] _T_1070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1786;
  reg [31:0] _T_1071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1787;
  reg [31:0] _T_1071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1788;
  reg [31:0] _T_1072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1789;
  reg [31:0] _T_1072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1790;
  reg [31:0] _T_1073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1791;
  reg [31:0] _T_1073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1792;
  reg [31:0] _T_1074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1793;
  reg [31:0] _T_1074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1794;
  reg [31:0] _T_1075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1795;
  reg [31:0] _T_1075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1796;
  reg [31:0] _T_1076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1797;
  reg [31:0] _T_1076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1798;
  reg [31:0] _T_1077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1799;
  reg [31:0] _T_1077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1800;
  reg [31:0] _T_1078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1801;
  reg [31:0] _T_1078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1802;
  reg [31:0] _T_1079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1803;
  reg [31:0] _T_1079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1804;
  reg [31:0] _T_1080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1805;
  reg [31:0] _T_1080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1806;
  reg [31:0] _T_1081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1807;
  reg [31:0] _T_1081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1808;
  reg [31:0] _T_1082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1809;
  reg [31:0] _T_1082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1810;
  reg [31:0] _T_1083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1811;
  reg [31:0] _T_1083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1812;
  reg [31:0] _T_1084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1813;
  reg [31:0] _T_1084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1814;
  reg [31:0] _T_1085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1815;
  reg [31:0] _T_1085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1816;
  reg [31:0] _T_1086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1817;
  reg [31:0] _T_1086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1818;
  reg [31:0] _T_1087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1819;
  reg [31:0] _T_1087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1820;
  reg [31:0] _T_1088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1821;
  reg [31:0] _T_1088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1822;
  reg [31:0] _T_1089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1823;
  reg [31:0] _T_1089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1824;
  reg [31:0] _T_1090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1825;
  reg [31:0] _T_1090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1826;
  reg [31:0] _T_1091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1827;
  reg [31:0] _T_1091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1828;
  reg [31:0] _T_1092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1829;
  reg [31:0] _T_1092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1830;
  reg [31:0] _T_1093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1831;
  reg [31:0] _T_1093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1832;
  reg [31:0] _T_1094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1833;
  reg [31:0] _T_1094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1834;
  reg [31:0] _T_1095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1835;
  reg [31:0] _T_1095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1836;
  reg [31:0] _T_1096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1837;
  reg [31:0] _T_1096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1838;
  reg [31:0] _T_1097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1839;
  reg [31:0] _T_1097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1840;
  reg [31:0] _T_1098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1841;
  reg [31:0] _T_1098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1842;
  reg [31:0] _T_1099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1843;
  reg [31:0] _T_1099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1844;
  reg [31:0] _T_1100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1845;
  reg [31:0] _T_1100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1846;
  reg [31:0] _T_1101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1847;
  reg [31:0] _T_1101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1848;
  reg [31:0] _T_1102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1849;
  reg [31:0] _T_1102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1850;
  reg [31:0] _T_1103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1851;
  reg [31:0] _T_1103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1852;
  reg [31:0] _T_1104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1853;
  reg [31:0] _T_1104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1854;
  reg [31:0] _T_1105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1855;
  reg [31:0] _T_1105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1856;
  reg [31:0] _T_1106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1857;
  reg [31:0] _T_1106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1858;
  reg [31:0] _T_1107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1859;
  reg [31:0] _T_1107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1860;
  reg [31:0] _T_1108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1861;
  reg [31:0] _T_1108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1862;
  reg [31:0] _T_1109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1863;
  reg [31:0] _T_1109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1864;
  reg [31:0] _T_1110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1865;
  reg [31:0] _T_1110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1866;
  reg [31:0] _T_1111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1867;
  reg [31:0] _T_1111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1868;
  reg [31:0] _T_1112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1869;
  reg [31:0] _T_1112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1870;
  reg [31:0] _T_1113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1871;
  reg [31:0] _T_1113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1872;
  reg [31:0] _T_1114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1873;
  reg [31:0] _T_1114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1874;
  reg [31:0] _T_1115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1875;
  reg [31:0] _T_1115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1876;
  reg [31:0] _T_1116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1877;
  reg [31:0] _T_1116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1878;
  reg [31:0] _T_1117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1879;
  reg [31:0] _T_1117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1880;
  reg [31:0] _T_1118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1881;
  reg [31:0] _T_1118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1882;
  reg [31:0] _T_1119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1883;
  reg [31:0] _T_1119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1884;
  reg [31:0] _T_1120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1885;
  reg [31:0] _T_1120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1886;
  reg [31:0] _T_1121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1887;
  reg [31:0] _T_1121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1888;
  reg [31:0] _T_1122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1889;
  reg [31:0] _T_1122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1890;
  reg [31:0] _T_1123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1891;
  reg [31:0] _T_1123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1892;
  reg [31:0] _T_1124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1893;
  reg [31:0] _T_1124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1894;
  reg [31:0] _T_1125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1895;
  reg [31:0] _T_1125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1896;
  reg [31:0] _T_1126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1897;
  reg [31:0] _T_1126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1898;
  reg [31:0] _T_1127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1899;
  reg [31:0] _T_1127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1900;
  reg [31:0] _T_1128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1901;
  reg [31:0] _T_1128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1902;
  reg [31:0] _T_1129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1903;
  reg [31:0] _T_1129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1904;
  reg [31:0] _T_1130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1905;
  reg [31:0] _T_1130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1906;
  reg [31:0] _T_1131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1907;
  reg [31:0] _T_1131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1908;
  reg [31:0] _T_1132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1909;
  reg [31:0] _T_1132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1910;
  reg [31:0] _T_1133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1911;
  reg [31:0] _T_1133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1912;
  reg [31:0] _T_1134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1913;
  reg [31:0] _T_1134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1914;
  reg [31:0] _T_1135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1915;
  reg [31:0] _T_1135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1916;
  reg [31:0] _T_1136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1917;
  reg [31:0] _T_1136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1918;
  reg [31:0] _T_1137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1919;
  reg [31:0] _T_1137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1920;
  reg [31:0] _T_1138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1921;
  reg [31:0] _T_1138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1922;
  reg [31:0] _T_1139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1923;
  reg [31:0] _T_1139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1924;
  reg [31:0] _T_1140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1925;
  reg [31:0] _T_1140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1926;
  reg [31:0] _T_1141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1927;
  reg [31:0] _T_1141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1928;
  reg [31:0] _T_1142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1929;
  reg [31:0] _T_1142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1930;
  reg [31:0] _T_1143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1931;
  reg [31:0] _T_1143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1932;
  reg [31:0] _T_1144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1933;
  reg [31:0] _T_1144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1934;
  reg [31:0] _T_1145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1935;
  reg [31:0] _T_1145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1936;
  reg [31:0] _T_1146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1937;
  reg [31:0] _T_1146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1938;
  reg [31:0] _T_1147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1939;
  reg [31:0] _T_1147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1940;
  reg [31:0] _T_1148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1941;
  reg [31:0] _T_1148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1942;
  reg [31:0] _T_1149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1943;
  reg [31:0] _T_1149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1944;
  reg [31:0] _T_1150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1945;
  reg [31:0] _T_1150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1946;
  reg [31:0] _T_1151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1947;
  reg [31:0] _T_1151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1948;
  reg [31:0] _T_1152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1949;
  reg [31:0] _T_1152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1950;
  reg [31:0] _T_1153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1951;
  reg [31:0] _T_1153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1952;
  reg [31:0] _T_1154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1953;
  reg [31:0] _T_1154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1954;
  reg [31:0] _T_1155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1955;
  reg [31:0] _T_1155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1956;
  reg [31:0] _T_1156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1957;
  reg [31:0] _T_1156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1958;
  reg [31:0] _T_1157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1959;
  reg [31:0] _T_1157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1960;
  reg [31:0] _T_1158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1961;
  reg [31:0] _T_1158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1962;
  reg [31:0] _T_1159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1963;
  reg [31:0] _T_1159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1964;
  reg [31:0] _T_1160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1965;
  reg [31:0] _T_1160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1966;
  reg [31:0] _T_1161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1967;
  reg [31:0] _T_1161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1968;
  reg [31:0] _T_1162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1969;
  reg [31:0] _T_1162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1970;
  reg [31:0] _T_1163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1971;
  reg [31:0] _T_1163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1972;
  reg [31:0] _T_1164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1973;
  reg [31:0] _T_1164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1974;
  reg [31:0] _T_1165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1975;
  reg [31:0] _T_1165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1976;
  reg [31:0] _T_1166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1977;
  reg [31:0] _T_1166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1978;
  reg [31:0] _T_1167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1979;
  reg [31:0] _T_1167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1980;
  reg [31:0] _T_1168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1981;
  reg [31:0] _T_1168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1982;
  reg [31:0] _T_1169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1983;
  reg [31:0] _T_1169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1984;
  reg [31:0] _T_1170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1985;
  reg [31:0] _T_1170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1986;
  reg [31:0] _T_1171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1987;
  reg [31:0] _T_1171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1988;
  reg [31:0] _T_1172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1989;
  reg [31:0] _T_1172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1990;
  reg [31:0] _T_1173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1991;
  reg [31:0] _T_1173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1992;
  reg [31:0] _T_1174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1993;
  reg [31:0] _T_1174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1994;
  reg [31:0] _T_1175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1995;
  reg [31:0] _T_1175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1996;
  reg [31:0] _T_1176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1997;
  reg [31:0] _T_1176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1998;
  reg [31:0] _T_1177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1999;
  reg [31:0] _T_1177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2000;
  reg [31:0] _T_1178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2001;
  reg [31:0] _T_1178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2002;
  reg [31:0] _T_1179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2003;
  reg [31:0] _T_1179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2004;
  reg [31:0] _T_1180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2005;
  reg [31:0] _T_1180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2006;
  reg [31:0] _T_1181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2007;
  reg [31:0] _T_1181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2008;
  reg [31:0] _T_1182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2009;
  reg [31:0] _T_1182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2010;
  reg [31:0] _T_1183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2011;
  reg [31:0] _T_1183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2012;
  reg [31:0] _T_1184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2013;
  reg [31:0] _T_1184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2014;
  reg [31:0] _T_1185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2015;
  reg [31:0] _T_1185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2016;
  reg [31:0] _T_1186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2017;
  reg [31:0] _T_1186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2018;
  reg [31:0] _T_1187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2019;
  reg [31:0] _T_1187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2020;
  reg [31:0] _T_1188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2021;
  reg [31:0] _T_1188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2022;
  reg [31:0] _T_1189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2023;
  reg [31:0] _T_1189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2024;
  reg [31:0] _T_1190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2025;
  reg [31:0] _T_1190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2026;
  reg [31:0] _T_1191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2027;
  reg [31:0] _T_1191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2028;
  reg [31:0] _T_1192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2029;
  reg [31:0] _T_1192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2030;
  reg [31:0] _T_1193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2031;
  reg [31:0] _T_1193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2032;
  reg [31:0] _T_1194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2033;
  reg [31:0] _T_1194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2034;
  reg [31:0] _T_1195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2035;
  reg [31:0] _T_1195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2036;
  reg [31:0] _T_1196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2037;
  reg [31:0] _T_1196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2038;
  reg [31:0] _T_1197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2039;
  reg [31:0] _T_1197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2040;
  reg [31:0] _T_1198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2041;
  reg [31:0] _T_1198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2042;
  reg [31:0] _T_1199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2043;
  reg [31:0] _T_1199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2044;
  reg [31:0] _T_1200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2045;
  reg [31:0] _T_1200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2046;
  reg [31:0] _T_1201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2047;
  reg [31:0] _T_1201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2048;
  reg [31:0] _T_1202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2049;
  reg [31:0] _T_1202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2050;
  reg [31:0] _T_1203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2051;
  reg [31:0] _T_1203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2052;
  reg [31:0] _T_1204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2053;
  reg [31:0] _T_1204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2054;
  reg [31:0] _T_1207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2055;
  reg [31:0] _T_1207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2056;
  reg [31:0] _T_1208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2057;
  reg [31:0] _T_1208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2058;
  reg [31:0] _T_1209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2059;
  reg [31:0] _T_1209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2060;
  reg [31:0] _T_1210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2061;
  reg [31:0] _T_1210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2062;
  reg [31:0] _T_1211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2063;
  reg [31:0] _T_1211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2064;
  reg [31:0] _T_1212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2065;
  reg [31:0] _T_1212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2066;
  reg [31:0] _T_1213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2067;
  reg [31:0] _T_1213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2068;
  reg [31:0] _T_1214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2069;
  reg [31:0] _T_1214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2070;
  reg [31:0] _T_1215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2071;
  reg [31:0] _T_1215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2072;
  reg [31:0] _T_1216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2073;
  reg [31:0] _T_1216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2074;
  reg [31:0] _T_1217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2075;
  reg [31:0] _T_1217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2076;
  reg [31:0] _T_1218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2077;
  reg [31:0] _T_1218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2078;
  reg [31:0] _T_1219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2079;
  reg [31:0] _T_1219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2080;
  reg [31:0] _T_1220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2081;
  reg [31:0] _T_1220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2082;
  reg [31:0] _T_1221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2083;
  reg [31:0] _T_1221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2084;
  reg [31:0] _T_1222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2085;
  reg [31:0] _T_1222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2086;
  reg [31:0] _T_1223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2087;
  reg [31:0] _T_1223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2088;
  reg [31:0] _T_1224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2089;
  reg [31:0] _T_1224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2090;
  reg [31:0] _T_1225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2091;
  reg [31:0] _T_1225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2092;
  reg [31:0] _T_1226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2093;
  reg [31:0] _T_1226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2094;
  reg [31:0] _T_1227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2095;
  reg [31:0] _T_1227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2096;
  reg [31:0] _T_1228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2097;
  reg [31:0] _T_1228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2098;
  reg [31:0] _T_1229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2099;
  reg [31:0] _T_1229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2100;
  reg [31:0] _T_1230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2101;
  reg [31:0] _T_1230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2102;
  reg [31:0] _T_1231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2103;
  reg [31:0] _T_1231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2104;
  reg [31:0] _T_1232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2105;
  reg [31:0] _T_1232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2106;
  reg [31:0] _T_1233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2107;
  reg [31:0] _T_1233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2108;
  reg [31:0] _T_1234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2109;
  reg [31:0] _T_1234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2110;
  reg [31:0] _T_1235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2111;
  reg [31:0] _T_1235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2112;
  reg [31:0] _T_1236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2113;
  reg [31:0] _T_1236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2114;
  reg [31:0] _T_1237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2115;
  reg [31:0] _T_1237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2116;
  reg [31:0] _T_1238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2117;
  reg [31:0] _T_1238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2118;
  reg [31:0] _T_1239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2119;
  reg [31:0] _T_1239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2120;
  reg [31:0] _T_1240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2121;
  reg [31:0] _T_1240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2122;
  reg [31:0] _T_1241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2123;
  reg [31:0] _T_1241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2124;
  reg [31:0] _T_1242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2125;
  reg [31:0] _T_1242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2126;
  reg [31:0] _T_1243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2127;
  reg [31:0] _T_1243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2128;
  reg [31:0] _T_1244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2129;
  reg [31:0] _T_1244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2130;
  reg [31:0] _T_1245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2131;
  reg [31:0] _T_1245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2132;
  reg [31:0] _T_1246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2133;
  reg [31:0] _T_1246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2134;
  reg [31:0] _T_1247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2135;
  reg [31:0] _T_1247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2136;
  reg [31:0] _T_1248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2137;
  reg [31:0] _T_1248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2138;
  reg [31:0] _T_1249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2139;
  reg [31:0] _T_1249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2140;
  reg [31:0] _T_1250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2141;
  reg [31:0] _T_1250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2142;
  reg [31:0] _T_1251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2143;
  reg [31:0] _T_1251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2144;
  reg [31:0] _T_1252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2145;
  reg [31:0] _T_1252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2146;
  reg [31:0] _T_1253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2147;
  reg [31:0] _T_1253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2148;
  reg [31:0] _T_1254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2149;
  reg [31:0] _T_1254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2150;
  reg [31:0] _T_1255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2151;
  reg [31:0] _T_1255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2152;
  reg [31:0] _T_1256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2153;
  reg [31:0] _T_1256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2154;
  reg [31:0] _T_1257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2155;
  reg [31:0] _T_1257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2156;
  reg [31:0] _T_1258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2157;
  reg [31:0] _T_1258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2158;
  reg [31:0] _T_1259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2159;
  reg [31:0] _T_1259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2160;
  reg [31:0] _T_1260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2161;
  reg [31:0] _T_1260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2162;
  reg [31:0] _T_1261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2163;
  reg [31:0] _T_1261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2164;
  reg [31:0] _T_1262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2165;
  reg [31:0] _T_1262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2166;
  reg [31:0] _T_1263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2167;
  reg [31:0] _T_1263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2168;
  reg [31:0] _T_1264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2169;
  reg [31:0] _T_1264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2170;
  reg [31:0] _T_1265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2171;
  reg [31:0] _T_1265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2172;
  reg [31:0] _T_1266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2173;
  reg [31:0] _T_1266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2174;
  reg [31:0] _T_1267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2175;
  reg [31:0] _T_1267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2176;
  reg [31:0] _T_1268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2177;
  reg [31:0] _T_1268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2178;
  reg [31:0] _T_1269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2179;
  reg [31:0] _T_1269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2180;
  reg [31:0] _T_1270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2181;
  reg [31:0] _T_1270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2182;
  reg [31:0] _T_1271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2183;
  reg [31:0] _T_1271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2184;
  reg [31:0] _T_1272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2185;
  reg [31:0] _T_1272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2186;
  reg [31:0] _T_1273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2187;
  reg [31:0] _T_1273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2188;
  reg [31:0] _T_1274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2189;
  reg [31:0] _T_1274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2190;
  reg [31:0] _T_1275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2191;
  reg [31:0] _T_1275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2192;
  reg [31:0] _T_1276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2193;
  reg [31:0] _T_1276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2194;
  reg [31:0] _T_1277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2195;
  reg [31:0] _T_1277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2196;
  reg [31:0] _T_1278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2197;
  reg [31:0] _T_1278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2198;
  reg [31:0] _T_1279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2199;
  reg [31:0] _T_1279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2200;
  reg [31:0] _T_1280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2201;
  reg [31:0] _T_1280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2202;
  reg [31:0] _T_1281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2203;
  reg [31:0] _T_1281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2204;
  reg [31:0] _T_1282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2205;
  reg [31:0] _T_1282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2206;
  reg [31:0] _T_1283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2207;
  reg [31:0] _T_1283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2208;
  reg [31:0] _T_1284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2209;
  reg [31:0] _T_1284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2210;
  reg [31:0] _T_1285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2211;
  reg [31:0] _T_1285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2212;
  reg [31:0] _T_1286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2213;
  reg [31:0] _T_1286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2214;
  reg [31:0] _T_1287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2215;
  reg [31:0] _T_1287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2216;
  reg [31:0] _T_1288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2217;
  reg [31:0] _T_1288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2218;
  reg [31:0] _T_1289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2219;
  reg [31:0] _T_1289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2220;
  reg [31:0] _T_1290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2221;
  reg [31:0] _T_1290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2222;
  reg [31:0] _T_1291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2223;
  reg [31:0] _T_1291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2224;
  reg [31:0] _T_1292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2225;
  reg [31:0] _T_1292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2226;
  reg [31:0] _T_1293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2227;
  reg [31:0] _T_1293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2228;
  reg [31:0] _T_1294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2229;
  reg [31:0] _T_1294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2230;
  reg [31:0] _T_1295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2231;
  reg [31:0] _T_1295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2232;
  reg [31:0] _T_1296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2233;
  reg [31:0] _T_1296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2234;
  reg [31:0] _T_1297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2235;
  reg [31:0] _T_1297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2236;
  reg [31:0] _T_1298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2237;
  reg [31:0] _T_1298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2238;
  reg [31:0] _T_1299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2239;
  reg [31:0] _T_1299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2240;
  reg [31:0] _T_1300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2241;
  reg [31:0] _T_1300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2242;
  reg [31:0] _T_1301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2243;
  reg [31:0] _T_1301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2244;
  reg [31:0] _T_1302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2245;
  reg [31:0] _T_1302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2246;
  reg [31:0] _T_1303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2247;
  reg [31:0] _T_1303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2248;
  reg [31:0] _T_1304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2249;
  reg [31:0] _T_1304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2250;
  reg [31:0] _T_1305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2251;
  reg [31:0] _T_1305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2252;
  reg [31:0] _T_1306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2253;
  reg [31:0] _T_1306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2254;
  reg [31:0] _T_1307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2255;
  reg [31:0] _T_1307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2256;
  reg [31:0] _T_1308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2257;
  reg [31:0] _T_1308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2258;
  reg [31:0] _T_1309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2259;
  reg [31:0] _T_1309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2260;
  reg [31:0] _T_1310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2261;
  reg [31:0] _T_1310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2262;
  reg [31:0] _T_1311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2263;
  reg [31:0] _T_1311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2264;
  reg [31:0] _T_1312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2265;
  reg [31:0] _T_1312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2266;
  reg [31:0] _T_1313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2267;
  reg [31:0] _T_1313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2268;
  reg [31:0] _T_1314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2269;
  reg [31:0] _T_1314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2270;
  reg [31:0] _T_1315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2271;
  reg [31:0] _T_1315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2272;
  reg [31:0] _T_1316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2273;
  reg [31:0] _T_1316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2274;
  reg [31:0] _T_1317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2275;
  reg [31:0] _T_1317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2276;
  reg [31:0] _T_1318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2277;
  reg [31:0] _T_1318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2278;
  reg [31:0] _T_1319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2279;
  reg [31:0] _T_1319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2280;
  reg [31:0] _T_1320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2281;
  reg [31:0] _T_1320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2282;
  reg [31:0] _T_1321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2283;
  reg [31:0] _T_1321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2284;
  reg [31:0] _T_1322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2285;
  reg [31:0] _T_1322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2286;
  reg [31:0] _T_1323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2287;
  reg [31:0] _T_1323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2288;
  reg [31:0] _T_1324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2289;
  reg [31:0] _T_1324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2290;
  reg [31:0] _T_1325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2291;
  reg [31:0] _T_1325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2292;
  reg [31:0] _T_1326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2293;
  reg [31:0] _T_1326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2294;
  reg [31:0] _T_1327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2295;
  reg [31:0] _T_1327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2296;
  reg [31:0] _T_1328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2297;
  reg [31:0] _T_1328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2298;
  reg [31:0] _T_1329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2299;
  reg [31:0] _T_1329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2300;
  reg [31:0] _T_1330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2301;
  reg [31:0] _T_1330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2302;
  reg [31:0] _T_1331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2303;
  reg [31:0] _T_1331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2304;
  reg [31:0] _T_1332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2305;
  reg [31:0] _T_1332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2306;
  reg [31:0] _T_1333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2307;
  reg [31:0] _T_1333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2308;
  reg [31:0] _T_1334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2309;
  reg [31:0] _T_1334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2310;
  reg [31:0] _T_1335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2311;
  reg [31:0] _T_1335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2312;
  reg [31:0] _T_1336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2313;
  reg [31:0] _T_1336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2314;
  reg [31:0] _T_1337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2315;
  reg [31:0] _T_1337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2316;
  reg [31:0] _T_1338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2317;
  reg [31:0] _T_1338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2318;
  reg [31:0] _T_1339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2319;
  reg [31:0] _T_1339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2320;
  reg [31:0] _T_1340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2321;
  reg [31:0] _T_1340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2322;
  reg [31:0] _T_1341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2323;
  reg [31:0] _T_1341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2324;
  reg [31:0] _T_1342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2325;
  reg [31:0] _T_1342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2326;
  reg [31:0] _T_1343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2327;
  reg [31:0] _T_1343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2328;
  reg [31:0] _T_1344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2329;
  reg [31:0] _T_1344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2330;
  reg [31:0] _T_1345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2331;
  reg [31:0] _T_1345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2332;
  reg [31:0] _T_1346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2333;
  reg [31:0] _T_1346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2334;
  reg [31:0] _T_1347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2335;
  reg [31:0] _T_1347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2336;
  reg [31:0] _T_1348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2337;
  reg [31:0] _T_1348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2338;
  reg [31:0] _T_1349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2339;
  reg [31:0] _T_1349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2340;
  reg [31:0] _T_1350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2341;
  reg [31:0] _T_1350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2342;
  reg [31:0] _T_1351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2343;
  reg [31:0] _T_1351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2344;
  reg [31:0] _T_1352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2345;
  reg [31:0] _T_1352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2346;
  reg [31:0] _T_1353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2347;
  reg [31:0] _T_1353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2348;
  reg [31:0] _T_1354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2349;
  reg [31:0] _T_1354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2350;
  reg [31:0] _T_1355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2351;
  reg [31:0] _T_1355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2352;
  reg [31:0] _T_1356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2353;
  reg [31:0] _T_1356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2354;
  reg [31:0] _T_1357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2355;
  reg [31:0] _T_1357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2356;
  reg [31:0] _T_1358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2357;
  reg [31:0] _T_1358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2358;
  reg [31:0] _T_1359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2359;
  reg [31:0] _T_1359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2360;
  reg [31:0] _T_1360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2361;
  reg [31:0] _T_1360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2362;
  reg [31:0] _T_1361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2363;
  reg [31:0] _T_1361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2364;
  reg [31:0] _T_1362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2365;
  reg [31:0] _T_1362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2366;
  reg [31:0] _T_1363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2367;
  reg [31:0] _T_1363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2368;
  reg [31:0] _T_1364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2369;
  reg [31:0] _T_1364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2370;
  reg [31:0] _T_1365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2371;
  reg [31:0] _T_1365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2372;
  reg [31:0] _T_1366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2373;
  reg [31:0] _T_1366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2374;
  reg [31:0] _T_1367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2375;
  reg [31:0] _T_1367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2376;
  reg [31:0] _T_1368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2377;
  reg [31:0] _T_1368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2378;
  reg [31:0] _T_1369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2379;
  reg [31:0] _T_1369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2380;
  reg [31:0] _T_1370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2381;
  reg [31:0] _T_1370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2382;
  reg [31:0] _T_1371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2383;
  reg [31:0] _T_1371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2384;
  reg [31:0] _T_1372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2385;
  reg [31:0] _T_1372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2386;
  reg [31:0] _T_1373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2387;
  reg [31:0] _T_1373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2388;
  reg [31:0] _T_1374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2389;
  reg [31:0] _T_1374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2390;
  reg [31:0] _T_1375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2391;
  reg [31:0] _T_1375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2392;
  reg [31:0] _T_1376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2393;
  reg [31:0] _T_1376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2394;
  reg [31:0] _T_1377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2395;
  reg [31:0] _T_1377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2396;
  reg [31:0] _T_1378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2397;
  reg [31:0] _T_1378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2398;
  reg [31:0] _T_1379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2399;
  reg [31:0] _T_1379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2400;
  reg [31:0] _T_1380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2401;
  reg [31:0] _T_1380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2402;
  reg [31:0] _T_1381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2403;
  reg [31:0] _T_1381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2404;
  reg [31:0] _T_1382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2405;
  reg [31:0] _T_1382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2406;
  reg [31:0] _T_1383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2407;
  reg [31:0] _T_1383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2408;
  reg [31:0] _T_1384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2409;
  reg [31:0] _T_1384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2410;
  reg [31:0] _T_1385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2411;
  reg [31:0] _T_1385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2412;
  reg [31:0] _T_1386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2413;
  reg [31:0] _T_1386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2414;
  reg [31:0] _T_1387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2415;
  reg [31:0] _T_1387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2416;
  reg [31:0] _T_1388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2417;
  reg [31:0] _T_1388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2418;
  reg [31:0] _T_1389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2419;
  reg [31:0] _T_1389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2420;
  reg [31:0] _T_1390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2421;
  reg [31:0] _T_1390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2422;
  reg [31:0] _T_1391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2423;
  reg [31:0] _T_1391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2424;
  reg [31:0] _T_1392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2425;
  reg [31:0] _T_1392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2426;
  reg [31:0] _T_1393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2427;
  reg [31:0] _T_1393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2428;
  reg [31:0] _T_1394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2429;
  reg [31:0] _T_1394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2430;
  reg [31:0] _T_1395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2431;
  reg [31:0] _T_1395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2432;
  reg [31:0] _T_1396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2433;
  reg [31:0] _T_1396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2434;
  reg [31:0] _T_1397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2435;
  reg [31:0] _T_1397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2436;
  reg [31:0] _T_1398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2437;
  reg [31:0] _T_1398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2438;
  reg [31:0] _T_1399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2439;
  reg [31:0] _T_1399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2440;
  reg [31:0] _T_1400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2441;
  reg [31:0] _T_1400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2442;
  reg [31:0] _T_1401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2443;
  reg [31:0] _T_1401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2444;
  reg [31:0] _T_1402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2445;
  reg [31:0] _T_1402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2446;
  reg [31:0] _T_1403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2447;
  reg [31:0] _T_1403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2448;
  reg [31:0] _T_1404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2449;
  reg [31:0] _T_1404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2450;
  reg [31:0] _T_1405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2451;
  reg [31:0] _T_1405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2452;
  reg [31:0] _T_1406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2453;
  reg [31:0] _T_1406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2454;
  reg [31:0] _T_1407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2455;
  reg [31:0] _T_1407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2456;
  reg [31:0] _T_1408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2457;
  reg [31:0] _T_1408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2458;
  reg [31:0] _T_1409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2459;
  reg [31:0] _T_1409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2460;
  reg [31:0] _T_1410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2461;
  reg [31:0] _T_1410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2462;
  reg [31:0] _T_1411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2463;
  reg [31:0] _T_1411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2464;
  reg [31:0] _T_1412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2465;
  reg [31:0] _T_1412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2466;
  reg [31:0] _T_1413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2467;
  reg [31:0] _T_1413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2468;
  reg [31:0] _T_1414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2469;
  reg [31:0] _T_1414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2470;
  reg [31:0] _T_1415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2471;
  reg [31:0] _T_1415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2472;
  reg [31:0] _T_1416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2473;
  reg [31:0] _T_1416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2474;
  reg [31:0] _T_1417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2475;
  reg [31:0] _T_1417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2476;
  reg [31:0] _T_1418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2477;
  reg [31:0] _T_1418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2478;
  reg [31:0] _T_1419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2479;
  reg [31:0] _T_1419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2480;
  reg [31:0] _T_1420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2481;
  reg [31:0] _T_1420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2482;
  reg [31:0] _T_1421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2483;
  reg [31:0] _T_1421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2484;
  reg [31:0] _T_1422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2485;
  reg [31:0] _T_1422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2486;
  reg [31:0] _T_1423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2487;
  reg [31:0] _T_1423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2488;
  reg [31:0] _T_1424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2489;
  reg [31:0] _T_1424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2490;
  reg [31:0] _T_1425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2491;
  reg [31:0] _T_1425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2492;
  reg [31:0] _T_1426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2493;
  reg [31:0] _T_1426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2494;
  reg [31:0] _T_1427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2495;
  reg [31:0] _T_1427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2496;
  reg [31:0] _T_1428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2497;
  reg [31:0] _T_1428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2498;
  reg [31:0] _T_1429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2499;
  reg [31:0] _T_1429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2500;
  reg [31:0] _T_1430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2501;
  reg [31:0] _T_1430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2502;
  reg [31:0] _T_1431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2503;
  reg [31:0] _T_1431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2504;
  reg [31:0] _T_1432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2505;
  reg [31:0] _T_1432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2506;
  reg [31:0] _T_1433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2507;
  reg [31:0] _T_1433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2508;
  reg [31:0] _T_1434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2509;
  reg [31:0] _T_1434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2510;
  reg [31:0] _T_1435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2511;
  reg [31:0] _T_1435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2512;
  reg [31:0] _T_1436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2513;
  reg [31:0] _T_1436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2514;
  reg [31:0] _T_1437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2515;
  reg [31:0] _T_1437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2516;
  reg [31:0] _T_1438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2517;
  reg [31:0] _T_1438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2518;
  reg [31:0] _T_1439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2519;
  reg [31:0] _T_1439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2520;
  reg [31:0] _T_1440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2521;
  reg [31:0] _T_1440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2522;
  reg [31:0] _T_1441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2523;
  reg [31:0] _T_1441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2524;
  reg [31:0] _T_1442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2525;
  reg [31:0] _T_1442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2526;
  reg [31:0] _T_1443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2527;
  reg [31:0] _T_1443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2528;
  reg [31:0] _T_1444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2529;
  reg [31:0] _T_1444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2530;
  reg [31:0] _T_1445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2531;
  reg [31:0] _T_1445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2532;
  reg [31:0] _T_1446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2533;
  reg [31:0] _T_1446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2534;
  reg [31:0] _T_1447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2535;
  reg [31:0] _T_1447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2536;
  reg [31:0] _T_1448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2537;
  reg [31:0] _T_1448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2538;
  reg [31:0] _T_1449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2539;
  reg [31:0] _T_1449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2540;
  reg [31:0] _T_1450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2541;
  reg [31:0] _T_1450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2542;
  reg [31:0] _T_1451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2543;
  reg [31:0] _T_1451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2544;
  reg [31:0] _T_1452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2545;
  reg [31:0] _T_1452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2546;
  reg [31:0] _T_1453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2547;
  reg [31:0] _T_1453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2548;
  reg [31:0] _T_1454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2549;
  reg [31:0] _T_1454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2550;
  reg [31:0] _T_1455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2551;
  reg [31:0] _T_1455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2552;
  reg [31:0] _T_1456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2553;
  reg [31:0] _T_1456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2554;
  reg [31:0] _T_1457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2555;
  reg [31:0] _T_1457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2556;
  reg [31:0] _T_1458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2557;
  reg [31:0] _T_1458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2558;
  reg [31:0] _T_1459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2559;
  reg [31:0] _T_1459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2560;
  reg [31:0] _T_1460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2561;
  reg [31:0] _T_1460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2562;
  reg [31:0] _T_1461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2563;
  reg [31:0] _T_1461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2564;
  reg [31:0] _T_1462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2565;
  reg [31:0] _T_1462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2566;
  reg [31:0] _T_1463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2567;
  reg [31:0] _T_1463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2568;
  reg [31:0] _T_1464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2569;
  reg [31:0] _T_1464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2570;
  reg [31:0] _T_1465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2571;
  reg [31:0] _T_1465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2572;
  reg [31:0] _T_1466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2573;
  reg [31:0] _T_1466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2574;
  reg [31:0] _T_1467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2575;
  reg [31:0] _T_1467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2576;
  reg [31:0] _T_1468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2577;
  reg [31:0] _T_1468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2578;
  reg [31:0] _T_1469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2579;
  reg [31:0] _T_1469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2580;
  reg [31:0] _T_1470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2581;
  reg [31:0] _T_1470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2582;
  reg [31:0] _T_1471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2583;
  reg [31:0] _T_1471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2584;
  reg [31:0] _T_1472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2585;
  reg [31:0] _T_1472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2586;
  reg [31:0] _T_1473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2587;
  reg [31:0] _T_1473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2588;
  reg [31:0] _T_1474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2589;
  reg [31:0] _T_1474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2590;
  reg [31:0] _T_1475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2591;
  reg [31:0] _T_1475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2592;
  reg [31:0] _T_1476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2593;
  reg [31:0] _T_1476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2594;
  reg [31:0] _T_1477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2595;
  reg [31:0] _T_1477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2596;
  reg [31:0] _T_1478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2597;
  reg [31:0] _T_1478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2598;
  reg [31:0] _T_1479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2599;
  reg [31:0] _T_1479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2600;
  reg [31:0] _T_1480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2601;
  reg [31:0] _T_1480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2602;
  reg [31:0] _T_1481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2603;
  reg [31:0] _T_1481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2604;
  reg [31:0] _T_1482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2605;
  reg [31:0] _T_1482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2606;
  reg [31:0] _T_1483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2607;
  reg [31:0] _T_1483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2608;
  reg [31:0] _T_1484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2609;
  reg [31:0] _T_1484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2610;
  reg [31:0] _T_1485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2611;
  reg [31:0] _T_1485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2612;
  reg [31:0] _T_1486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2613;
  reg [31:0] _T_1486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2614;
  reg [31:0] _T_1487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2615;
  reg [31:0] _T_1487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2616;
  reg [31:0] _T_1488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2617;
  reg [31:0] _T_1488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2618;
  reg [31:0] _T_1489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2619;
  reg [31:0] _T_1489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2620;
  reg [31:0] _T_1490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2621;
  reg [31:0] _T_1490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2622;
  reg [31:0] _T_1491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2623;
  reg [31:0] _T_1491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2624;
  reg [31:0] _T_1492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2625;
  reg [31:0] _T_1492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2626;
  reg [31:0] _T_1493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2627;
  reg [31:0] _T_1493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2628;
  reg [31:0] _T_1494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2629;
  reg [31:0] _T_1494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2630;
  reg [31:0] _T_1495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2631;
  reg [31:0] _T_1495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2632;
  reg [31:0] _T_1496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2633;
  reg [31:0] _T_1496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2634;
  reg [31:0] _T_1497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2635;
  reg [31:0] _T_1497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2636;
  reg [31:0] _T_1498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2637;
  reg [31:0] _T_1498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2638;
  reg [31:0] _T_1499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2639;
  reg [31:0] _T_1499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2640;
  reg [31:0] _T_1500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2641;
  reg [31:0] _T_1500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2642;
  reg [31:0] _T_1501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2643;
  reg [31:0] _T_1501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2644;
  reg [31:0] _T_1502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2645;
  reg [31:0] _T_1502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2646;
  reg [31:0] _T_1503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2647;
  reg [31:0] _T_1503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2648;
  reg [31:0] _T_1504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2649;
  reg [31:0] _T_1504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2650;
  reg [31:0] _T_1505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2651;
  reg [31:0] _T_1505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2652;
  reg [31:0] _T_1506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2653;
  reg [31:0] _T_1506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2654;
  reg [31:0] _T_1507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2655;
  reg [31:0] _T_1507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2656;
  reg [31:0] _T_1508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2657;
  reg [31:0] _T_1508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2658;
  reg [31:0] _T_1509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2659;
  reg [31:0] _T_1509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2660;
  reg [31:0] _T_1510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2661;
  reg [31:0] _T_1510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2662;
  reg [31:0] _T_1511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2663;
  reg [31:0] _T_1511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2664;
  reg [31:0] _T_1512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2665;
  reg [31:0] _T_1512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2666;
  reg [31:0] _T_1513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2667;
  reg [31:0] _T_1513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2668;
  reg [31:0] _T_1514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2669;
  reg [31:0] _T_1514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2670;
  reg [31:0] _T_1515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2671;
  reg [31:0] _T_1515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2672;
  reg [31:0] _T_1516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2673;
  reg [31:0] _T_1516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2674;
  reg [31:0] _T_1517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2675;
  reg [31:0] _T_1517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2676;
  reg [31:0] _T_1518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2677;
  reg [31:0] _T_1518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2678;
  reg [31:0] _T_1519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2679;
  reg [31:0] _T_1519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2680;
  reg [31:0] _T_1520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2681;
  reg [31:0] _T_1520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2682;
  reg [31:0] _T_1521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2683;
  reg [31:0] _T_1521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2684;
  reg [31:0] _T_1522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2685;
  reg [31:0] _T_1522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2686;
  reg [31:0] _T_1523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2687;
  reg [31:0] _T_1523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2688;
  reg [31:0] _T_1524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2689;
  reg [31:0] _T_1524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2690;
  reg [31:0] _T_1525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2691;
  reg [31:0] _T_1525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2692;
  reg [31:0] _T_1526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2693;
  reg [31:0] _T_1526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2694;
  reg [31:0] _T_1527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2695;
  reg [31:0] _T_1527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2696;
  reg [31:0] _T_1528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2697;
  reg [31:0] _T_1528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2698;
  reg [31:0] _T_1529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2699;
  reg [31:0] _T_1529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2700;
  reg [31:0] _T_1530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2701;
  reg [31:0] _T_1530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2702;
  reg [31:0] _T_1531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2703;
  reg [31:0] _T_1531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2704;
  reg [31:0] _T_1532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2705;
  reg [31:0] _T_1532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2706;
  reg [31:0] _T_1533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2707;
  reg [31:0] _T_1533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2708;
  reg [31:0] _T_1534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2709;
  reg [31:0] _T_1534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2710;
  reg [31:0] _T_1535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2711;
  reg [31:0] _T_1535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2712;
  reg [31:0] _T_1536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2713;
  reg [31:0] _T_1536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2714;
  reg [31:0] _T_1537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2715;
  reg [31:0] _T_1537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2716;
  reg [31:0] _T_1538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2717;
  reg [31:0] _T_1538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2718;
  reg [31:0] _T_1539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2719;
  reg [31:0] _T_1539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2720;
  reg [31:0] _T_1540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2721;
  reg [31:0] _T_1540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2722;
  reg [31:0] _T_1541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2723;
  reg [31:0] _T_1541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2724;
  reg [31:0] _T_1542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2725;
  reg [31:0] _T_1542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2726;
  reg [31:0] _T_1543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2727;
  reg [31:0] _T_1543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2728;
  reg [31:0] _T_1544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2729;
  reg [31:0] _T_1544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2730;
  reg [31:0] _T_1545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2731;
  reg [31:0] _T_1545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2732;
  reg [31:0] _T_1546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2733;
  reg [31:0] _T_1546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2734;
  reg [31:0] _T_1547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2735;
  reg [31:0] _T_1547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2736;
  reg [31:0] _T_1548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2737;
  reg [31:0] _T_1548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2738;
  reg [31:0] _T_1549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2739;
  reg [31:0] _T_1549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2740;
  reg [31:0] _T_1550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2741;
  reg [31:0] _T_1550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2742;
  reg [31:0] _T_1551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2743;
  reg [31:0] _T_1551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2744;
  reg [31:0] _T_1552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2745;
  reg [31:0] _T_1552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2746;
  reg [31:0] _T_1553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2747;
  reg [31:0] _T_1553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2748;
  reg [31:0] _T_1554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2749;
  reg [31:0] _T_1554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2750;
  reg [31:0] _T_1555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2751;
  reg [31:0] _T_1555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2752;
  reg [31:0] _T_1556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2753;
  reg [31:0] _T_1556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2754;
  reg [31:0] _T_1557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2755;
  reg [31:0] _T_1557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2756;
  reg [31:0] _T_1558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2757;
  reg [31:0] _T_1558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2758;
  reg [31:0] _T_1559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2759;
  reg [31:0] _T_1559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2760;
  reg [31:0] _T_1560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2761;
  reg [31:0] _T_1560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2762;
  reg [31:0] _T_1561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2763;
  reg [31:0] _T_1561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2764;
  reg [31:0] _T_1562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2765;
  reg [31:0] _T_1562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2766;
  reg [31:0] _T_1563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2767;
  reg [31:0] _T_1563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2768;
  reg [31:0] _T_1564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2769;
  reg [31:0] _T_1564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2770;
  reg [31:0] _T_1565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2771;
  reg [31:0] _T_1565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2772;
  reg [31:0] _T_1566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2773;
  reg [31:0] _T_1566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2774;
  reg [31:0] _T_1567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2775;
  reg [31:0] _T_1567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2776;
  reg [31:0] _T_1568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2777;
  reg [31:0] _T_1568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2778;
  reg [31:0] _T_1569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2779;
  reg [31:0] _T_1569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2780;
  reg [31:0] _T_1570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2781;
  reg [31:0] _T_1570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2782;
  reg [31:0] _T_1571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2783;
  reg [31:0] _T_1571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2784;
  reg [31:0] _T_1572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2785;
  reg [31:0] _T_1572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2786;
  reg [31:0] _T_1573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2787;
  reg [31:0] _T_1573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2788;
  reg [31:0] _T_1574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2789;
  reg [31:0] _T_1574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2790;
  reg [31:0] _T_1575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2791;
  reg [31:0] _T_1575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2792;
  reg [31:0] _T_1576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2793;
  reg [31:0] _T_1576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2794;
  reg [31:0] _T_1577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2795;
  reg [31:0] _T_1577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2796;
  reg [31:0] _T_1578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2797;
  reg [31:0] _T_1578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2798;
  reg [31:0] _T_1579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2799;
  reg [31:0] _T_1579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2800;
  reg [31:0] _T_1580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2801;
  reg [31:0] _T_1580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2802;
  reg [31:0] _T_1581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2803;
  reg [31:0] _T_1581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2804;
  reg [31:0] _T_1582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2805;
  reg [31:0] _T_1582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2806;
  reg [31:0] _T_1583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2807;
  reg [31:0] _T_1583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2808;
  reg [31:0] _T_1584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2809;
  reg [31:0] _T_1584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2810;
  reg [31:0] _T_1585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2811;
  reg [31:0] _T_1585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2812;
  reg [31:0] _T_1586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2813;
  reg [31:0] _T_1586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2814;
  reg [31:0] _T_1587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2815;
  reg [31:0] _T_1587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2816;
  reg [31:0] _T_1588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2817;
  reg [31:0] _T_1588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2818;
  reg [31:0] _T_1589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2819;
  reg [31:0] _T_1589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2820;
  reg [31:0] _T_1590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2821;
  reg [31:0] _T_1590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2822;
  reg [31:0] _T_1591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2823;
  reg [31:0] _T_1591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2824;
  reg [31:0] _T_1592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2825;
  reg [31:0] _T_1592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2826;
  reg [31:0] _T_1593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2827;
  reg [31:0] _T_1593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2828;
  reg [31:0] _T_1594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2829;
  reg [31:0] _T_1594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2830;
  reg [31:0] _T_1595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2831;
  reg [31:0] _T_1595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2832;
  reg [31:0] _T_1596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2833;
  reg [31:0] _T_1596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2834;
  reg [31:0] _T_1597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2835;
  reg [31:0] _T_1597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2836;
  reg [31:0] _T_1598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2837;
  reg [31:0] _T_1598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2838;
  reg [31:0] _T_1599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2839;
  reg [31:0] _T_1599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2840;
  reg [31:0] _T_1600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2841;
  reg [31:0] _T_1600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2842;
  reg [31:0] _T_1601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2843;
  reg [31:0] _T_1601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2844;
  reg [31:0] _T_1602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2845;
  reg [31:0] _T_1602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2846;
  reg [31:0] _T_1603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2847;
  reg [31:0] _T_1603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2848;
  reg [31:0] _T_1604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2849;
  reg [31:0] _T_1604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2850;
  reg [31:0] _T_1605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2851;
  reg [31:0] _T_1605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2852;
  reg [31:0] _T_1606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2853;
  reg [31:0] _T_1606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2854;
  reg [31:0] _T_1607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2855;
  reg [31:0] _T_1607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2856;
  reg [31:0] _T_1608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2857;
  reg [31:0] _T_1608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2858;
  reg [31:0] _T_1609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2859;
  reg [31:0] _T_1609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2860;
  reg [31:0] _T_1610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2861;
  reg [31:0] _T_1610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2862;
  reg [31:0] _T_1611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2863;
  reg [31:0] _T_1611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2864;
  reg [31:0] _T_1612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2865;
  reg [31:0] _T_1612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2866;
  reg [31:0] _T_1613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2867;
  reg [31:0] _T_1613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2868;
  reg [31:0] _T_1614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2869;
  reg [31:0] _T_1614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2870;
  reg [31:0] _T_1615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2871;
  reg [31:0] _T_1615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2872;
  reg [31:0] _T_1616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2873;
  reg [31:0] _T_1616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2874;
  reg [31:0] _T_1617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2875;
  reg [31:0] _T_1617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2876;
  reg [31:0] _T_1618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2877;
  reg [31:0] _T_1618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2878;
  reg [31:0] _T_1619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2879;
  reg [31:0] _T_1619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2880;
  reg [31:0] _T_1620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2881;
  reg [31:0] _T_1620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2882;
  reg [31:0] _T_1621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2883;
  reg [31:0] _T_1621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2884;
  reg [31:0] _T_1622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2885;
  reg [31:0] _T_1622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2886;
  reg [31:0] _T_1623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2887;
  reg [31:0] _T_1623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2888;
  reg [31:0] _T_1624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2889;
  reg [31:0] _T_1624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2890;
  reg [31:0] _T_1625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2891;
  reg [31:0] _T_1625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2892;
  reg [31:0] _T_1626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2893;
  reg [31:0] _T_1626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2894;
  reg [31:0] _T_1627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2895;
  reg [31:0] _T_1627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2896;
  reg [31:0] _T_1628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2897;
  reg [31:0] _T_1628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2898;
  reg [31:0] _T_1629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2899;
  reg [31:0] _T_1629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2900;
  reg [31:0] _T_1630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2901;
  reg [31:0] _T_1630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2902;
  reg [31:0] _T_1631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2903;
  reg [31:0] _T_1631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2904;
  reg [31:0] _T_1632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2905;
  reg [31:0] _T_1632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2906;
  reg [31:0] _T_1633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2907;
  reg [31:0] _T_1633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2908;
  reg [31:0] _T_1634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2909;
  reg [31:0] _T_1634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2910;
  reg [31:0] _T_1635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2911;
  reg [31:0] _T_1635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2912;
  reg [31:0] _T_1636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2913;
  reg [31:0] _T_1636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2914;
  reg [31:0] _T_1637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2915;
  reg [31:0] _T_1637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2916;
  reg [31:0] _T_1638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2917;
  reg [31:0] _T_1638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2918;
  reg [31:0] _T_1639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2919;
  reg [31:0] _T_1639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2920;
  reg [31:0] _T_1640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2921;
  reg [31:0] _T_1640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2922;
  reg [31:0] _T_1641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2923;
  reg [31:0] _T_1641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2924;
  reg [31:0] _T_1642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2925;
  reg [31:0] _T_1642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2926;
  reg [31:0] _T_1643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2927;
  reg [31:0] _T_1643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2928;
  reg [31:0] _T_1644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2929;
  reg [31:0] _T_1644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2930;
  reg [31:0] _T_1645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2931;
  reg [31:0] _T_1645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2932;
  reg [31:0] _T_1646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2933;
  reg [31:0] _T_1646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2934;
  reg [31:0] _T_1647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2935;
  reg [31:0] _T_1647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2936;
  reg [31:0] _T_1648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2937;
  reg [31:0] _T_1648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2938;
  reg [31:0] _T_1649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2939;
  reg [31:0] _T_1649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2940;
  reg [31:0] _T_1650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2941;
  reg [31:0] _T_1650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2942;
  reg [31:0] _T_1651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2943;
  reg [31:0] _T_1651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2944;
  reg [31:0] _T_1652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2945;
  reg [31:0] _T_1652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2946;
  reg [31:0] _T_1653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2947;
  reg [31:0] _T_1653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2948;
  reg [31:0] _T_1654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2949;
  reg [31:0] _T_1654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2950;
  reg [31:0] _T_1655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2951;
  reg [31:0] _T_1655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2952;
  reg [31:0] _T_1656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2953;
  reg [31:0] _T_1656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2954;
  reg [31:0] _T_1657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2955;
  reg [31:0] _T_1657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2956;
  reg [31:0] _T_1658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2957;
  reg [31:0] _T_1658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2958;
  reg [31:0] _T_1659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2959;
  reg [31:0] _T_1659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2960;
  reg [31:0] _T_1660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2961;
  reg [31:0] _T_1660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2962;
  reg [31:0] _T_1661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2963;
  reg [31:0] _T_1661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2964;
  reg [31:0] _T_1662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2965;
  reg [31:0] _T_1662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2966;
  reg [31:0] _T_1663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2967;
  reg [31:0] _T_1663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2968;
  reg [31:0] _T_1664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2969;
  reg [31:0] _T_1664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2970;
  reg [31:0] _T_1665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2971;
  reg [31:0] _T_1665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2972;
  reg [31:0] _T_1666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2973;
  reg [31:0] _T_1666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2974;
  reg [31:0] _T_1667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2975;
  reg [31:0] _T_1667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2976;
  reg [31:0] _T_1668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2977;
  reg [31:0] _T_1668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2978;
  reg [31:0] _T_1669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2979;
  reg [31:0] _T_1669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2980;
  reg [31:0] _T_1670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2981;
  reg [31:0] _T_1670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2982;
  reg [31:0] _T_1671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2983;
  reg [31:0] _T_1671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2984;
  reg [31:0] _T_1672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2985;
  reg [31:0] _T_1672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2986;
  reg [31:0] _T_1673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2987;
  reg [31:0] _T_1673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2988;
  reg [31:0] _T_1674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2989;
  reg [31:0] _T_1674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2990;
  reg [31:0] _T_1675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2991;
  reg [31:0] _T_1675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2992;
  reg [31:0] _T_1676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2993;
  reg [31:0] _T_1676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2994;
  reg [31:0] _T_1677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2995;
  reg [31:0] _T_1677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2996;
  reg [31:0] _T_1678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2997;
  reg [31:0] _T_1678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2998;
  reg [31:0] _T_1679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2999;
  reg [31:0] _T_1679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3000;
  reg [31:0] _T_1680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3001;
  reg [31:0] _T_1680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3002;
  reg [31:0] _T_1681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3003;
  reg [31:0] _T_1681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3004;
  reg [31:0] _T_1682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3005;
  reg [31:0] _T_1682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3006;
  reg [31:0] _T_1683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3007;
  reg [31:0] _T_1683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3008;
  reg [31:0] _T_1684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3009;
  reg [31:0] _T_1684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3010;
  reg [31:0] _T_1685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3011;
  reg [31:0] _T_1685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3012;
  reg [31:0] _T_1686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3013;
  reg [31:0] _T_1686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3014;
  reg [31:0] _T_1687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3015;
  reg [31:0] _T_1687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3016;
  reg [31:0] _T_1688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3017;
  reg [31:0] _T_1688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3018;
  reg [31:0] _T_1689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3019;
  reg [31:0] _T_1689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3020;
  reg [31:0] _T_1690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3021;
  reg [31:0] _T_1690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3022;
  reg [31:0] _T_1691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3023;
  reg [31:0] _T_1691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3024;
  reg [31:0] _T_1692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3025;
  reg [31:0] _T_1692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3026;
  reg [31:0] _T_1693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3027;
  reg [31:0] _T_1693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3028;
  reg [31:0] _T_1694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3029;
  reg [31:0] _T_1694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3030;
  reg [31:0] _T_1695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3031;
  reg [31:0] _T_1695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3032;
  reg [31:0] _T_1696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3033;
  reg [31:0] _T_1696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3034;
  reg [31:0] _T_1697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3035;
  reg [31:0] _T_1697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3036;
  reg [31:0] _T_1698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3037;
  reg [31:0] _T_1698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3038;
  reg [31:0] _T_1699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3039;
  reg [31:0] _T_1699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3040;
  reg [31:0] _T_1700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3041;
  reg [31:0] _T_1700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3042;
  reg [31:0] _T_1701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3043;
  reg [31:0] _T_1701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3044;
  reg [31:0] _T_1702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3045;
  reg [31:0] _T_1702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3046;
  reg [31:0] _T_1703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3047;
  reg [31:0] _T_1703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3048;
  reg [31:0] _T_1704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3049;
  reg [31:0] _T_1704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3050;
  reg [31:0] _T_1705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3051;
  reg [31:0] _T_1705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3052;
  reg [31:0] _T_1706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3053;
  reg [31:0] _T_1706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3054;
  reg [31:0] _T_1707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3055;
  reg [31:0] _T_1707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3056;
  reg [31:0] _T_1708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3057;
  reg [31:0] _T_1708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3058;
  reg [31:0] _T_1709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3059;
  reg [31:0] _T_1709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3060;
  reg [31:0] _T_1710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3061;
  reg [31:0] _T_1710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3062;
  reg [31:0] _T_1711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3063;
  reg [31:0] _T_1711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3064;
  reg [31:0] _T_1712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3065;
  reg [31:0] _T_1712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3066;
  reg [31:0] _T_1713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3067;
  reg [31:0] _T_1713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3068;
  reg [31:0] _T_1714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3069;
  reg [31:0] _T_1714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3070;
  reg [31:0] _T_1715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3071;
  reg [31:0] _T_1715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3072;
  reg [31:0] _T_1716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3073;
  reg [31:0] _T_1716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3074;
  reg [31:0] _T_1717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3075;
  reg [31:0] _T_1717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3076;
  reg [31:0] _T_1718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3077;
  reg [31:0] _T_1718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3078;
  wire [63:0] _T_1723;
  reg [31:0] _T_1728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3079;
  reg [31:0] _T_1728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3080;
  reg [31:0] _T_1729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3081;
  reg [31:0] _T_1729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3082;
  reg [31:0] _T_1730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3083;
  reg [31:0] _T_1730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3084;
  reg [31:0] _T_1731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3085;
  reg [31:0] _T_1731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3086;
  reg [31:0] _T_1732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3087;
  reg [31:0] _T_1732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3088;
  reg [31:0] _T_1733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3089;
  reg [31:0] _T_1733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3090;
  reg [31:0] _T_1734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3091;
  reg [31:0] _T_1734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3092;
  reg [31:0] _T_1735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3093;
  reg [31:0] _T_1735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3094;
  reg [31:0] _T_1736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3095;
  reg [31:0] _T_1736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3096;
  reg [31:0] _T_1737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3097;
  reg [31:0] _T_1737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3098;
  reg [31:0] _T_1738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3099;
  reg [31:0] _T_1738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3100;
  reg [31:0] _T_1739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3101;
  reg [31:0] _T_1739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3102;
  reg [31:0] _T_1740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3103;
  reg [31:0] _T_1740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3104;
  reg [31:0] _T_1741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3105;
  reg [31:0] _T_1741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3106;
  reg [31:0] _T_1742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3107;
  reg [31:0] _T_1742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3108;
  reg [31:0] _T_1743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3109;
  reg [31:0] _T_1743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3110;
  reg [31:0] _T_1744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3111;
  reg [31:0] _T_1744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3112;
  reg [31:0] _T_1745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3113;
  reg [31:0] _T_1745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3114;
  reg [31:0] _T_1746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3115;
  reg [31:0] _T_1746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3116;
  reg [31:0] _T_1747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3117;
  reg [31:0] _T_1747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3118;
  reg [31:0] _T_1748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3119;
  reg [31:0] _T_1748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3120;
  reg [31:0] _T_1749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3121;
  reg [31:0] _T_1749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3122;
  reg [31:0] _T_1750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3123;
  reg [31:0] _T_1750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3124;
  reg [31:0] _T_1751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3125;
  reg [31:0] _T_1751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3126;
  reg [31:0] _T_1752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3127;
  reg [31:0] _T_1752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3128;
  reg [31:0] _T_1753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3129;
  reg [31:0] _T_1753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3130;
  reg [31:0] _T_1754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3131;
  reg [31:0] _T_1754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3132;
  reg [31:0] _T_1755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3133;
  reg [31:0] _T_1755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3134;
  reg [31:0] _T_1756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3135;
  reg [31:0] _T_1756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3136;
  reg [31:0] _T_1757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3137;
  reg [31:0] _T_1757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3138;
  reg [31:0] _T_1758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3139;
  reg [31:0] _T_1758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3140;
  reg [31:0] _T_1759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3141;
  reg [31:0] _T_1759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3142;
  reg [31:0] _T_1760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3143;
  reg [31:0] _T_1760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3144;
  reg [31:0] _T_1761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3145;
  reg [31:0] _T_1761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3146;
  reg [31:0] _T_1762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3147;
  reg [31:0] _T_1762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3148;
  reg [31:0] _T_1763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3149;
  reg [31:0] _T_1763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3150;
  reg [31:0] _T_1764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3151;
  reg [31:0] _T_1764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3152;
  reg [31:0] _T_1765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3153;
  reg [31:0] _T_1765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3154;
  reg [31:0] _T_1766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3155;
  reg [31:0] _T_1766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3156;
  reg [31:0] _T_1767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3157;
  reg [31:0] _T_1767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3158;
  reg [31:0] _T_1768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3159;
  reg [31:0] _T_1768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3160;
  reg [31:0] _T_1769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3161;
  reg [31:0] _T_1769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3162;
  reg [31:0] _T_1770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3163;
  reg [31:0] _T_1770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3164;
  reg [31:0] _T_1771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3165;
  reg [31:0] _T_1771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3166;
  reg [31:0] _T_1772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3167;
  reg [31:0] _T_1772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3168;
  reg [31:0] _T_1773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3169;
  reg [31:0] _T_1773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3170;
  reg [31:0] _T_1774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3171;
  reg [31:0] _T_1774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3172;
  reg [31:0] _T_1775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3173;
  reg [31:0] _T_1775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3174;
  reg [31:0] _T_1776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3175;
  reg [31:0] _T_1776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3176;
  reg [31:0] _T_1777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3177;
  reg [31:0] _T_1777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3178;
  reg [31:0] _T_1778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3179;
  reg [31:0] _T_1778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3180;
  reg [31:0] _T_1779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3181;
  reg [31:0] _T_1779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3182;
  reg [31:0] _T_1780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3183;
  reg [31:0] _T_1780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3184;
  reg [31:0] _T_1781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3185;
  reg [31:0] _T_1781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3186;
  reg [31:0] _T_1782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3187;
  reg [31:0] _T_1782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3188;
  reg [31:0] _T_1783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3189;
  reg [31:0] _T_1783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3190;
  reg [31:0] _T_1784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3191;
  reg [31:0] _T_1784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3192;
  reg [31:0] _T_1785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3193;
  reg [31:0] _T_1785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3194;
  reg [31:0] _T_1786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3195;
  reg [31:0] _T_1786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3196;
  reg [31:0] _T_1787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3197;
  reg [31:0] _T_1787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3198;
  reg [31:0] _T_1788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3199;
  reg [31:0] _T_1788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3200;
  reg [31:0] _T_1789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3201;
  reg [31:0] _T_1789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3202;
  reg [31:0] _T_1790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3203;
  reg [31:0] _T_1790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3204;
  reg [31:0] _T_1791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3205;
  reg [31:0] _T_1791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3206;
  reg [31:0] _T_1792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3207;
  reg [31:0] _T_1792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3208;
  reg [31:0] _T_1793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3209;
  reg [31:0] _T_1793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3210;
  reg [31:0] _T_1794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3211;
  reg [31:0] _T_1794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3212;
  reg [31:0] _T_1795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3213;
  reg [31:0] _T_1795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3214;
  reg [31:0] _T_1796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3215;
  reg [31:0] _T_1796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3216;
  reg [31:0] _T_1797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3217;
  reg [31:0] _T_1797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3218;
  reg [31:0] _T_1798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3219;
  reg [31:0] _T_1798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3220;
  reg [31:0] _T_1799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3221;
  reg [31:0] _T_1799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3222;
  reg [31:0] _T_1800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3223;
  reg [31:0] _T_1800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3224;
  reg [31:0] _T_1801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3225;
  reg [31:0] _T_1801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3226;
  reg [31:0] _T_1802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3227;
  reg [31:0] _T_1802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3228;
  reg [31:0] _T_1803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3229;
  reg [31:0] _T_1803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3230;
  reg [31:0] _T_1804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3231;
  reg [31:0] _T_1804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3232;
  reg [31:0] _T_1805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3233;
  reg [31:0] _T_1805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3234;
  reg [31:0] _T_1806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3235;
  reg [31:0] _T_1806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3236;
  reg [31:0] _T_1807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3237;
  reg [31:0] _T_1807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3238;
  reg [31:0] _T_1808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3239;
  reg [31:0] _T_1808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3240;
  reg [31:0] _T_1809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3241;
  reg [31:0] _T_1809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3242;
  reg [31:0] _T_1810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3243;
  reg [31:0] _T_1810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3244;
  reg [31:0] _T_1811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3245;
  reg [31:0] _T_1811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3246;
  reg [31:0] _T_1812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3247;
  reg [31:0] _T_1812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3248;
  reg [31:0] _T_1813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3249;
  reg [31:0] _T_1813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3250;
  reg [31:0] _T_1814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3251;
  reg [31:0] _T_1814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3252;
  reg [31:0] _T_1815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3253;
  reg [31:0] _T_1815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3254;
  reg [31:0] _T_1816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3255;
  reg [31:0] _T_1816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3256;
  reg [31:0] _T_1817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3257;
  reg [31:0] _T_1817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3258;
  reg [31:0] _T_1818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3259;
  reg [31:0] _T_1818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3260;
  reg [31:0] _T_1819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3261;
  reg [31:0] _T_1819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3262;
  reg [31:0] _T_1820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3263;
  reg [31:0] _T_1820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3264;
  reg [31:0] _T_1821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3265;
  reg [31:0] _T_1821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3266;
  reg [31:0] _T_1822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3267;
  reg [31:0] _T_1822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3268;
  reg [31:0] _T_1823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3269;
  reg [31:0] _T_1823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3270;
  reg [31:0] _T_1824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3271;
  reg [31:0] _T_1824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3272;
  reg [31:0] _T_1825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3273;
  reg [31:0] _T_1825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3274;
  reg [31:0] _T_1826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3275;
  reg [31:0] _T_1826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3276;
  reg [31:0] _T_1827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3277;
  reg [31:0] _T_1827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3278;
  reg [31:0] _T_1828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3279;
  reg [31:0] _T_1828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3280;
  reg [31:0] _T_1829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3281;
  reg [31:0] _T_1829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3282;
  reg [31:0] _T_1830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3283;
  reg [31:0] _T_1830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3284;
  reg [31:0] _T_1831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3285;
  reg [31:0] _T_1831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3286;
  reg [31:0] _T_1832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3287;
  reg [31:0] _T_1832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3288;
  reg [31:0] _T_1833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3289;
  reg [31:0] _T_1833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3290;
  reg [31:0] _T_1834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3291;
  reg [31:0] _T_1834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3292;
  reg [31:0] _T_1835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3293;
  reg [31:0] _T_1835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3294;
  reg [31:0] _T_1836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3295;
  reg [31:0] _T_1836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3296;
  reg [31:0] _T_1837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3297;
  reg [31:0] _T_1837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3298;
  reg [31:0] _T_1838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3299;
  reg [31:0] _T_1838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3300;
  reg [31:0] _T_1839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3301;
  reg [31:0] _T_1839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3302;
  reg [31:0] _T_1840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3303;
  reg [31:0] _T_1840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3304;
  reg [31:0] _T_1841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3305;
  reg [31:0] _T_1841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3306;
  reg [31:0] _T_1842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3307;
  reg [31:0] _T_1842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3308;
  reg [31:0] _T_1843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3309;
  reg [31:0] _T_1843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3310;
  reg [31:0] _T_1844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3311;
  reg [31:0] _T_1844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3312;
  reg [31:0] _T_1845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3313;
  reg [31:0] _T_1845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3314;
  reg [31:0] _T_1846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3315;
  reg [31:0] _T_1846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3316;
  reg [31:0] _T_1847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3317;
  reg [31:0] _T_1847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3318;
  reg [31:0] _T_1848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3319;
  reg [31:0] _T_1848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3320;
  reg [31:0] _T_1849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3321;
  reg [31:0] _T_1849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3322;
  reg [31:0] _T_1850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3323;
  reg [31:0] _T_1850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3324;
  reg [31:0] _T_1851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3325;
  reg [31:0] _T_1851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3326;
  reg [31:0] _T_1852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3327;
  reg [31:0] _T_1852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3328;
  reg [31:0] _T_1853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3329;
  reg [31:0] _T_1853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3330;
  reg [31:0] _T_1854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3331;
  reg [31:0] _T_1854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3332;
  reg [31:0] _T_1855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3333;
  reg [31:0] _T_1855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3334;
  reg [31:0] _T_1856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3335;
  reg [31:0] _T_1856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3336;
  reg [31:0] _T_1857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3337;
  reg [31:0] _T_1857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3338;
  reg [31:0] _T_1858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3339;
  reg [31:0] _T_1858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3340;
  reg [31:0] _T_1859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3341;
  reg [31:0] _T_1859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3342;
  reg [31:0] _T_1860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3343;
  reg [31:0] _T_1860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3344;
  reg [31:0] _T_1861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3345;
  reg [31:0] _T_1861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3346;
  reg [31:0] _T_1862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3347;
  reg [31:0] _T_1862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3348;
  reg [31:0] _T_1863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3349;
  reg [31:0] _T_1863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3350;
  reg [31:0] _T_1864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3351;
  reg [31:0] _T_1864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3352;
  reg [31:0] _T_1865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3353;
  reg [31:0] _T_1865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3354;
  reg [31:0] _T_1866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3355;
  reg [31:0] _T_1866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3356;
  reg [31:0] _T_1867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3357;
  reg [31:0] _T_1867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3358;
  reg [31:0] _T_1868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3359;
  reg [31:0] _T_1868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3360;
  reg [31:0] _T_1869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3361;
  reg [31:0] _T_1869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3362;
  reg [31:0] _T_1870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3363;
  reg [31:0] _T_1870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3364;
  reg [31:0] _T_1871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3365;
  reg [31:0] _T_1871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3366;
  reg [31:0] _T_1872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3367;
  reg [31:0] _T_1872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3368;
  reg [31:0] _T_1873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3369;
  reg [31:0] _T_1873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3370;
  reg [31:0] _T_1874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3371;
  reg [31:0] _T_1874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3372;
  reg [31:0] _T_1875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3373;
  reg [31:0] _T_1875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3374;
  reg [31:0] _T_1876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3375;
  reg [31:0] _T_1876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3376;
  reg [31:0] _T_1877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3377;
  reg [31:0] _T_1877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3378;
  reg [31:0] _T_1878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3379;
  reg [31:0] _T_1878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3380;
  reg [31:0] _T_1879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3381;
  reg [31:0] _T_1879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3382;
  reg [31:0] _T_1880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3383;
  reg [31:0] _T_1880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3384;
  reg [31:0] _T_1881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3385;
  reg [31:0] _T_1881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3386;
  reg [31:0] _T_1882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3387;
  reg [31:0] _T_1882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3388;
  reg [31:0] _T_1883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3389;
  reg [31:0] _T_1883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3390;
  reg [31:0] _T_1884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3391;
  reg [31:0] _T_1884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3392;
  reg [31:0] _T_1885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3393;
  reg [31:0] _T_1885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3394;
  reg [31:0] _T_1886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3395;
  reg [31:0] _T_1886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3396;
  reg [31:0] _T_1887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3397;
  reg [31:0] _T_1887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3398;
  reg [31:0] _T_1888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3399;
  reg [31:0] _T_1888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3400;
  reg [31:0] _T_1889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3401;
  reg [31:0] _T_1889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3402;
  reg [31:0] _T_1890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3403;
  reg [31:0] _T_1890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3404;
  reg [31:0] _T_1891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3405;
  reg [31:0] _T_1891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3406;
  reg [31:0] _T_1892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3407;
  reg [31:0] _T_1892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3408;
  reg [31:0] _T_1893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3409;
  reg [31:0] _T_1893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3410;
  reg [31:0] _T_1894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3411;
  reg [31:0] _T_1894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3412;
  reg [31:0] _T_1895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3413;
  reg [31:0] _T_1895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3414;
  reg [31:0] _T_1896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3415;
  reg [31:0] _T_1896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3416;
  reg [31:0] _T_1897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3417;
  reg [31:0] _T_1897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3418;
  reg [31:0] _T_1898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3419;
  reg [31:0] _T_1898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3420;
  reg [31:0] _T_1899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3421;
  reg [31:0] _T_1899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3422;
  reg [31:0] _T_1900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3423;
  reg [31:0] _T_1900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3424;
  reg [31:0] _T_1901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3425;
  reg [31:0] _T_1901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3426;
  reg [31:0] _T_1902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3427;
  reg [31:0] _T_1902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3428;
  reg [31:0] _T_1903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3429;
  reg [31:0] _T_1903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3430;
  reg [31:0] _T_1904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3431;
  reg [31:0] _T_1904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3432;
  reg [31:0] _T_1905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3433;
  reg [31:0] _T_1905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3434;
  reg [31:0] _T_1906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3435;
  reg [31:0] _T_1906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3436;
  reg [31:0] _T_1907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3437;
  reg [31:0] _T_1907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3438;
  reg [31:0] _T_1908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3439;
  reg [31:0] _T_1908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3440;
  reg [31:0] _T_1909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3441;
  reg [31:0] _T_1909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3442;
  reg [31:0] _T_1910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3443;
  reg [31:0] _T_1910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3444;
  reg [31:0] _T_1911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3445;
  reg [31:0] _T_1911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3446;
  reg [31:0] _T_1912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3447;
  reg [31:0] _T_1912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3448;
  reg [31:0] _T_1913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3449;
  reg [31:0] _T_1913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3450;
  reg [31:0] _T_1914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3451;
  reg [31:0] _T_1914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3452;
  reg [31:0] _T_1915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3453;
  reg [31:0] _T_1915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3454;
  reg [31:0] _T_1916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3455;
  reg [31:0] _T_1916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3456;
  reg [31:0] _T_1917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3457;
  reg [31:0] _T_1917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3458;
  reg [31:0] _T_1918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3459;
  reg [31:0] _T_1918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3460;
  reg [31:0] _T_1919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3461;
  reg [31:0] _T_1919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3462;
  reg [31:0] _T_1920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3463;
  reg [31:0] _T_1920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3464;
  reg [31:0] _T_1921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3465;
  reg [31:0] _T_1921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3466;
  reg [31:0] _T_1922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3467;
  reg [31:0] _T_1922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3468;
  reg [31:0] _T_1923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3469;
  reg [31:0] _T_1923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3470;
  reg [31:0] _T_1924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3471;
  reg [31:0] _T_1924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3472;
  reg [31:0] _T_1925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3473;
  reg [31:0] _T_1925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3474;
  reg [31:0] _T_1926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3475;
  reg [31:0] _T_1926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3476;
  reg [31:0] _T_1927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3477;
  reg [31:0] _T_1927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3478;
  reg [31:0] _T_1928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3479;
  reg [31:0] _T_1928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3480;
  reg [31:0] _T_1929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3481;
  reg [31:0] _T_1929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3482;
  reg [31:0] _T_1930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3483;
  reg [31:0] _T_1930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3484;
  reg [31:0] _T_1931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3485;
  reg [31:0] _T_1931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3486;
  reg [31:0] _T_1932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3487;
  reg [31:0] _T_1932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3488;
  reg [31:0] _T_1933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3489;
  reg [31:0] _T_1933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3490;
  reg [31:0] _T_1934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3491;
  reg [31:0] _T_1934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3492;
  reg [31:0] _T_1935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3493;
  reg [31:0] _T_1935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3494;
  reg [31:0] _T_1936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3495;
  reg [31:0] _T_1936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3496;
  reg [31:0] _T_1937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3497;
  reg [31:0] _T_1937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3498;
  reg [31:0] _T_1938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3499;
  reg [31:0] _T_1938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3500;
  reg [31:0] _T_1939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3501;
  reg [31:0] _T_1939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3502;
  reg [31:0] _T_1940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3503;
  reg [31:0] _T_1940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3504;
  reg [31:0] _T_1941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3505;
  reg [31:0] _T_1941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3506;
  reg [31:0] _T_1942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3507;
  reg [31:0] _T_1942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3508;
  reg [31:0] _T_1943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3509;
  reg [31:0] _T_1943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3510;
  reg [31:0] _T_1944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3511;
  reg [31:0] _T_1944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3512;
  reg [31:0] _T_1945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3513;
  reg [31:0] _T_1945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3514;
  reg [31:0] _T_1946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3515;
  reg [31:0] _T_1946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3516;
  reg [31:0] _T_1947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3517;
  reg [31:0] _T_1947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3518;
  reg [31:0] _T_1948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3519;
  reg [31:0] _T_1948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3520;
  reg [31:0] _T_1949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3521;
  reg [31:0] _T_1949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3522;
  reg [31:0] _T_1950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3523;
  reg [31:0] _T_1950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3524;
  reg [31:0] _T_1951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3525;
  reg [31:0] _T_1951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3526;
  reg [31:0] _T_1952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3527;
  reg [31:0] _T_1952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3528;
  reg [31:0] _T_1953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3529;
  reg [31:0] _T_1953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3530;
  reg [31:0] _T_1954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3531;
  reg [31:0] _T_1954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3532;
  reg [31:0] _T_1955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3533;
  reg [31:0] _T_1955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3534;
  reg [31:0] _T_1956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3535;
  reg [31:0] _T_1956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3536;
  reg [31:0] _T_1957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3537;
  reg [31:0] _T_1957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3538;
  reg [31:0] _T_1958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3539;
  reg [31:0] _T_1958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3540;
  reg [31:0] _T_1959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3541;
  reg [31:0] _T_1959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3542;
  reg [31:0] _T_1960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3543;
  reg [31:0] _T_1960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3544;
  reg [31:0] _T_1961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3545;
  reg [31:0] _T_1961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3546;
  reg [31:0] _T_1962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3547;
  reg [31:0] _T_1962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3548;
  reg [31:0] _T_1963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3549;
  reg [31:0] _T_1963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3550;
  reg [31:0] _T_1964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3551;
  reg [31:0] _T_1964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3552;
  reg [31:0] _T_1965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3553;
  reg [31:0] _T_1965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3554;
  reg [31:0] _T_1966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3555;
  reg [31:0] _T_1966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3556;
  reg [31:0] _T_1967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3557;
  reg [31:0] _T_1967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3558;
  reg [31:0] _T_1968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3559;
  reg [31:0] _T_1968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3560;
  reg [31:0] _T_1969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3561;
  reg [31:0] _T_1969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3562;
  reg [31:0] _T_1970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3563;
  reg [31:0] _T_1970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3564;
  reg [31:0] _T_1971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3565;
  reg [31:0] _T_1971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3566;
  reg [31:0] _T_1972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3567;
  reg [31:0] _T_1972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3568;
  reg [31:0] _T_1973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3569;
  reg [31:0] _T_1973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3570;
  reg [31:0] _T_1974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3571;
  reg [31:0] _T_1974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3572;
  reg [31:0] _T_1975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3573;
  reg [31:0] _T_1975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3574;
  reg [31:0] _T_1976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3575;
  reg [31:0] _T_1976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3576;
  reg [31:0] _T_1977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3577;
  reg [31:0] _T_1977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3578;
  reg [31:0] _T_1978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3579;
  reg [31:0] _T_1978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3580;
  reg [31:0] _T_1979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3581;
  reg [31:0] _T_1979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3582;
  reg [31:0] _T_1980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3583;
  reg [31:0] _T_1980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3584;
  reg [31:0] _T_1981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3585;
  reg [31:0] _T_1981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3586;
  reg [31:0] _T_1982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3587;
  reg [31:0] _T_1982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3588;
  reg [31:0] _T_1983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3589;
  reg [31:0] _T_1983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3590;
  reg [31:0] _T_1984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3591;
  reg [31:0] _T_1984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3592;
  reg [31:0] _T_1985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3593;
  reg [31:0] _T_1985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3594;
  reg [31:0] _T_1986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3595;
  reg [31:0] _T_1986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3596;
  reg [31:0] _T_1987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3597;
  reg [31:0] _T_1987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3598;
  reg [31:0] _T_1988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3599;
  reg [31:0] _T_1988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3600;
  reg [31:0] _T_1989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3601;
  reg [31:0] _T_1989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3602;
  reg [31:0] _T_1990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3603;
  reg [31:0] _T_1990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3604;
  reg [31:0] _T_1991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3605;
  reg [31:0] _T_1991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3606;
  reg [31:0] _T_1992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3607;
  reg [31:0] _T_1992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3608;
  reg [31:0] _T_1993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3609;
  reg [31:0] _T_1993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3610;
  reg [31:0] _T_1994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3611;
  reg [31:0] _T_1994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3612;
  reg [31:0] _T_1995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3613;
  reg [31:0] _T_1995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3614;
  reg [31:0] _T_1996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3615;
  reg [31:0] _T_1996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3616;
  reg [31:0] _T_1997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3617;
  reg [31:0] _T_1997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3618;
  reg [31:0] _T_1998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3619;
  reg [31:0] _T_1998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3620;
  reg [31:0] _T_1999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3621;
  reg [31:0] _T_1999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3622;
  reg [31:0] _T_2000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3623;
  reg [31:0] _T_2000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3624;
  reg [31:0] _T_2001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3625;
  reg [31:0] _T_2001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3626;
  reg [31:0] _T_2002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3627;
  reg [31:0] _T_2002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3628;
  reg [31:0] _T_2003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3629;
  reg [31:0] _T_2003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3630;
  reg [31:0] _T_2004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3631;
  reg [31:0] _T_2004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3632;
  reg [31:0] _T_2005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3633;
  reg [31:0] _T_2005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3634;
  reg [31:0] _T_2006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3635;
  reg [31:0] _T_2006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3636;
  reg [31:0] _T_2007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3637;
  reg [31:0] _T_2007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3638;
  reg [31:0] _T_2008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3639;
  reg [31:0] _T_2008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3640;
  reg [31:0] _T_2009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3641;
  reg [31:0] _T_2009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3642;
  reg [31:0] _T_2010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3643;
  reg [31:0] _T_2010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3644;
  reg [31:0] _T_2011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3645;
  reg [31:0] _T_2011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3646;
  reg [31:0] _T_2012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3647;
  reg [31:0] _T_2012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3648;
  reg [31:0] _T_2013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3649;
  reg [31:0] _T_2013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3650;
  reg [31:0] _T_2014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3651;
  reg [31:0] _T_2014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3652;
  reg [31:0] _T_2015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3653;
  reg [31:0] _T_2015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3654;
  reg [31:0] _T_2016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3655;
  reg [31:0] _T_2016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3656;
  reg [31:0] _T_2017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3657;
  reg [31:0] _T_2017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3658;
  reg [31:0] _T_2018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3659;
  reg [31:0] _T_2018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3660;
  reg [31:0] _T_2019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3661;
  reg [31:0] _T_2019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3662;
  reg [31:0] _T_2020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3663;
  reg [31:0] _T_2020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3664;
  reg [31:0] _T_2021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3665;
  reg [31:0] _T_2021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3666;
  reg [31:0] _T_2022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3667;
  reg [31:0] _T_2022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3668;
  reg [31:0] _T_2023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3669;
  reg [31:0] _T_2023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3670;
  reg [31:0] _T_2024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3671;
  reg [31:0] _T_2024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3672;
  reg [31:0] _T_2025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3673;
  reg [31:0] _T_2025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3674;
  reg [31:0] _T_2026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3675;
  reg [31:0] _T_2026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3676;
  reg [31:0] _T_2027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3677;
  reg [31:0] _T_2027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3678;
  reg [31:0] _T_2028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3679;
  reg [31:0] _T_2028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3680;
  reg [31:0] _T_2029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3681;
  reg [31:0] _T_2029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3682;
  reg [31:0] _T_2030_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3683;
  reg [31:0] _T_2030_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3684;
  reg [31:0] _T_2031_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3685;
  reg [31:0] _T_2031_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3686;
  reg [31:0] _T_2032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3687;
  reg [31:0] _T_2032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3688;
  reg [31:0] _T_2033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3689;
  reg [31:0] _T_2033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3690;
  reg [31:0] _T_2034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3691;
  reg [31:0] _T_2034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3692;
  reg [31:0] _T_2035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3693;
  reg [31:0] _T_2035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3694;
  reg [31:0] _T_2036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3695;
  reg [31:0] _T_2036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3696;
  reg [31:0] _T_2037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3697;
  reg [31:0] _T_2037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3698;
  reg [31:0] _T_2038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3699;
  reg [31:0] _T_2038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3700;
  reg [31:0] _T_2039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3701;
  reg [31:0] _T_2039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3702;
  reg [31:0] _T_2040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3703;
  reg [31:0] _T_2040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3704;
  reg [31:0] _T_2041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3705;
  reg [31:0] _T_2041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3706;
  reg [31:0] _T_2042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3707;
  reg [31:0] _T_2042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3708;
  reg [31:0] _T_2043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3709;
  reg [31:0] _T_2043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3710;
  reg [31:0] _T_2044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3711;
  reg [31:0] _T_2044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3712;
  reg [31:0] _T_2045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3713;
  reg [31:0] _T_2045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3714;
  reg [31:0] _T_2046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3715;
  reg [31:0] _T_2046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3716;
  reg [31:0] _T_2047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3717;
  reg [31:0] _T_2047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3718;
  reg [31:0] _T_2048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3719;
  reg [31:0] _T_2048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3720;
  reg [31:0] _T_2049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3721;
  reg [31:0] _T_2049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3722;
  reg [31:0] _T_2050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3723;
  reg [31:0] _T_2050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3724;
  reg [31:0] _T_2051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3725;
  reg [31:0] _T_2051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3726;
  reg [31:0] _T_2052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3727;
  reg [31:0] _T_2052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3728;
  reg [31:0] _T_2053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3729;
  reg [31:0] _T_2053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3730;
  reg [31:0] _T_2054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3731;
  reg [31:0] _T_2054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3732;
  reg [31:0] _T_2055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3733;
  reg [31:0] _T_2055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3734;
  reg [31:0] _T_2056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3735;
  reg [31:0] _T_2056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3736;
  reg [31:0] _T_2057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3737;
  reg [31:0] _T_2057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3738;
  reg [31:0] _T_2058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3739;
  reg [31:0] _T_2058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3740;
  reg [31:0] _T_2059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3741;
  reg [31:0] _T_2059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3742;
  reg [31:0] _T_2060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3743;
  reg [31:0] _T_2060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3744;
  reg [31:0] _T_2061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3745;
  reg [31:0] _T_2061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3746;
  reg [31:0] _T_2062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3747;
  reg [31:0] _T_2062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3748;
  reg [31:0] _T_2063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3749;
  reg [31:0] _T_2063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3750;
  reg [31:0] _T_2064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3751;
  reg [31:0] _T_2064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3752;
  reg [31:0] _T_2065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3753;
  reg [31:0] _T_2065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3754;
  reg [31:0] _T_2066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3755;
  reg [31:0] _T_2066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3756;
  reg [31:0] _T_2067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3757;
  reg [31:0] _T_2067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3758;
  reg [31:0] _T_2068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3759;
  reg [31:0] _T_2068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3760;
  reg [31:0] _T_2069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3761;
  reg [31:0] _T_2069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3762;
  reg [31:0] _T_2070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3763;
  reg [31:0] _T_2070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3764;
  reg [31:0] _T_2071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3765;
  reg [31:0] _T_2071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3766;
  reg [31:0] _T_2072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3767;
  reg [31:0] _T_2072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3768;
  reg [31:0] _T_2073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3769;
  reg [31:0] _T_2073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3770;
  reg [31:0] _T_2074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3771;
  reg [31:0] _T_2074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3772;
  reg [31:0] _T_2075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3773;
  reg [31:0] _T_2075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3774;
  reg [31:0] _T_2076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3775;
  reg [31:0] _T_2076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3776;
  reg [31:0] _T_2077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3777;
  reg [31:0] _T_2077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3778;
  reg [31:0] _T_2078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3779;
  reg [31:0] _T_2078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3780;
  reg [31:0] _T_2079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3781;
  reg [31:0] _T_2079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3782;
  reg [31:0] _T_2080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3783;
  reg [31:0] _T_2080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3784;
  reg [31:0] _T_2081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3785;
  reg [31:0] _T_2081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3786;
  reg [31:0] _T_2082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3787;
  reg [31:0] _T_2082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3788;
  reg [31:0] _T_2083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3789;
  reg [31:0] _T_2083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3790;
  reg [31:0] _T_2084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3791;
  reg [31:0] _T_2084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3792;
  reg [31:0] _T_2085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3793;
  reg [31:0] _T_2085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3794;
  reg [31:0] _T_2086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3795;
  reg [31:0] _T_2086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3796;
  reg [31:0] _T_2087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3797;
  reg [31:0] _T_2087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3798;
  reg [31:0] _T_2088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3799;
  reg [31:0] _T_2088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3800;
  reg [31:0] _T_2089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3801;
  reg [31:0] _T_2089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3802;
  reg [31:0] _T_2090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3803;
  reg [31:0] _T_2090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3804;
  reg [31:0] _T_2091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3805;
  reg [31:0] _T_2091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3806;
  reg [31:0] _T_2092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3807;
  reg [31:0] _T_2092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3808;
  reg [31:0] _T_2093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3809;
  reg [31:0] _T_2093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3810;
  reg [31:0] _T_2094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3811;
  reg [31:0] _T_2094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3812;
  reg [31:0] _T_2095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3813;
  reg [31:0] _T_2095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3814;
  reg [31:0] _T_2096_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3815;
  reg [31:0] _T_2096_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3816;
  reg [31:0] _T_2097_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3817;
  reg [31:0] _T_2097_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3818;
  reg [31:0] _T_2098_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3819;
  reg [31:0] _T_2098_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3820;
  reg [31:0] _T_2099_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3821;
  reg [31:0] _T_2099_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3822;
  reg [31:0] _T_2100_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3823;
  reg [31:0] _T_2100_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3824;
  reg [31:0] _T_2101_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3825;
  reg [31:0] _T_2101_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3826;
  reg [31:0] _T_2102_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3827;
  reg [31:0] _T_2102_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3828;
  reg [31:0] _T_2103_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3829;
  reg [31:0] _T_2103_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3830;
  reg [31:0] _T_2104_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3831;
  reg [31:0] _T_2104_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3832;
  reg [31:0] _T_2105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3833;
  reg [31:0] _T_2105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3834;
  reg [31:0] _T_2106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3835;
  reg [31:0] _T_2106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3836;
  reg [31:0] _T_2107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3837;
  reg [31:0] _T_2107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3838;
  reg [31:0] _T_2108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3839;
  reg [31:0] _T_2108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3840;
  reg [31:0] _T_2109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3841;
  reg [31:0] _T_2109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3842;
  reg [31:0] _T_2110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3843;
  reg [31:0] _T_2110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3844;
  reg [31:0] _T_2111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3845;
  reg [31:0] _T_2111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3846;
  reg [31:0] _T_2112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3847;
  reg [31:0] _T_2112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3848;
  reg [31:0] _T_2113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3849;
  reg [31:0] _T_2113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3850;
  reg [31:0] _T_2114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3851;
  reg [31:0] _T_2114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3852;
  reg [31:0] _T_2115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3853;
  reg [31:0] _T_2115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3854;
  reg [31:0] _T_2116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3855;
  reg [31:0] _T_2116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3856;
  reg [31:0] _T_2117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3857;
  reg [31:0] _T_2117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3858;
  reg [31:0] _T_2118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3859;
  reg [31:0] _T_2118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3860;
  reg [31:0] _T_2119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3861;
  reg [31:0] _T_2119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3862;
  reg [31:0] _T_2120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3863;
  reg [31:0] _T_2120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3864;
  reg [31:0] _T_2121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3865;
  reg [31:0] _T_2121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3866;
  reg [31:0] _T_2122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3867;
  reg [31:0] _T_2122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3868;
  reg [31:0] _T_2123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3869;
  reg [31:0] _T_2123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3870;
  reg [31:0] _T_2124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3871;
  reg [31:0] _T_2124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3872;
  reg [31:0] _T_2125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3873;
  reg [31:0] _T_2125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3874;
  reg [31:0] _T_2126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3875;
  reg [31:0] _T_2126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3876;
  reg [31:0] _T_2127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3877;
  reg [31:0] _T_2127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3878;
  reg [31:0] _T_2128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3879;
  reg [31:0] _T_2128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3880;
  reg [31:0] _T_2129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3881;
  reg [31:0] _T_2129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3882;
  reg [31:0] _T_2130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3883;
  reg [31:0] _T_2130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3884;
  reg [31:0] _T_2131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3885;
  reg [31:0] _T_2131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3886;
  reg [31:0] _T_2132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3887;
  reg [31:0] _T_2132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3888;
  reg [31:0] _T_2133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3889;
  reg [31:0] _T_2133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3890;
  reg [31:0] _T_2134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3891;
  reg [31:0] _T_2134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3892;
  reg [31:0] _T_2135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3893;
  reg [31:0] _T_2135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3894;
  reg [31:0] _T_2136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3895;
  reg [31:0] _T_2136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3896;
  reg [31:0] _T_2137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3897;
  reg [31:0] _T_2137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3898;
  reg [31:0] _T_2138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3899;
  reg [31:0] _T_2138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3900;
  reg [31:0] _T_2139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3901;
  reg [31:0] _T_2139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3902;
  reg [31:0] _T_2140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3903;
  reg [31:0] _T_2140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3904;
  reg [31:0] _T_2141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3905;
  reg [31:0] _T_2141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3906;
  reg [31:0] _T_2142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3907;
  reg [31:0] _T_2142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3908;
  reg [31:0] _T_2143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3909;
  reg [31:0] _T_2143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3910;
  reg [31:0] _T_2144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3911;
  reg [31:0] _T_2144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3912;
  reg [31:0] _T_2145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3913;
  reg [31:0] _T_2145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3914;
  reg [31:0] _T_2146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3915;
  reg [31:0] _T_2146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3916;
  reg [31:0] _T_2147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3917;
  reg [31:0] _T_2147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3918;
  reg [31:0] _T_2148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3919;
  reg [31:0] _T_2148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3920;
  reg [31:0] _T_2149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3921;
  reg [31:0] _T_2149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3922;
  reg [31:0] _T_2150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3923;
  reg [31:0] _T_2150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3924;
  reg [31:0] _T_2151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3925;
  reg [31:0] _T_2151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3926;
  reg [31:0] _T_2152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3927;
  reg [31:0] _T_2152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3928;
  reg [31:0] _T_2153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3929;
  reg [31:0] _T_2153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3930;
  reg [31:0] _T_2154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3931;
  reg [31:0] _T_2154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3932;
  reg [31:0] _T_2155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3933;
  reg [31:0] _T_2155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3934;
  reg [31:0] _T_2156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3935;
  reg [31:0] _T_2156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3936;
  reg [31:0] _T_2157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3937;
  reg [31:0] _T_2157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3938;
  reg [31:0] _T_2158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3939;
  reg [31:0] _T_2158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3940;
  reg [31:0] _T_2159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3941;
  reg [31:0] _T_2159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3942;
  reg [31:0] _T_2160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3943;
  reg [31:0] _T_2160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3944;
  reg [31:0] _T_2161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3945;
  reg [31:0] _T_2161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3946;
  reg [31:0] _T_2162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3947;
  reg [31:0] _T_2162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3948;
  reg [31:0] _T_2163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3949;
  reg [31:0] _T_2163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3950;
  reg [31:0] _T_2164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3951;
  reg [31:0] _T_2164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3952;
  reg [31:0] _T_2165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3953;
  reg [31:0] _T_2165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3954;
  reg [31:0] _T_2166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3955;
  reg [31:0] _T_2166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3956;
  reg [31:0] _T_2167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3957;
  reg [31:0] _T_2167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3958;
  reg [31:0] _T_2168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3959;
  reg [31:0] _T_2168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3960;
  reg [31:0] _T_2169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3961;
  reg [31:0] _T_2169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3962;
  reg [31:0] _T_2170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3963;
  reg [31:0] _T_2170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3964;
  reg [31:0] _T_2171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3965;
  reg [31:0] _T_2171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3966;
  reg [31:0] _T_2172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3967;
  reg [31:0] _T_2172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3968;
  reg [31:0] _T_2173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3969;
  reg [31:0] _T_2173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3970;
  reg [31:0] _T_2174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3971;
  reg [31:0] _T_2174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3972;
  reg [31:0] _T_2175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3973;
  reg [31:0] _T_2175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3974;
  reg [31:0] _T_2176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3975;
  reg [31:0] _T_2176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3976;
  reg [31:0] _T_2177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3977;
  reg [31:0] _T_2177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3978;
  reg [31:0] _T_2178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3979;
  reg [31:0] _T_2178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3980;
  reg [31:0] _T_2179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3981;
  reg [31:0] _T_2179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3982;
  reg [31:0] _T_2180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3983;
  reg [31:0] _T_2180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3984;
  reg [31:0] _T_2181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3985;
  reg [31:0] _T_2181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3986;
  reg [31:0] _T_2182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3987;
  reg [31:0] _T_2182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3988;
  reg [31:0] _T_2183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3989;
  reg [31:0] _T_2183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3990;
  reg [31:0] _T_2184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3991;
  reg [31:0] _T_2184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3992;
  reg [31:0] _T_2185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3993;
  reg [31:0] _T_2185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3994;
  reg [31:0] _T_2186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3995;
  reg [31:0] _T_2186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3996;
  reg [31:0] _T_2187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3997;
  reg [31:0] _T_2187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3998;
  reg [31:0] _T_2188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3999;
  reg [31:0] _T_2188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4000;
  reg [31:0] _T_2189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4001;
  reg [31:0] _T_2189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4002;
  reg [31:0] _T_2190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4003;
  reg [31:0] _T_2190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4004;
  reg [31:0] _T_2191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4005;
  reg [31:0] _T_2191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4006;
  reg [31:0] _T_2192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4007;
  reg [31:0] _T_2192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4008;
  reg [31:0] _T_2193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4009;
  reg [31:0] _T_2193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4010;
  reg [31:0] _T_2194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4011;
  reg [31:0] _T_2194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4012;
  reg [31:0] _T_2195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4013;
  reg [31:0] _T_2195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4014;
  reg [31:0] _T_2196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4015;
  reg [31:0] _T_2196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4016;
  reg [31:0] _T_2197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4017;
  reg [31:0] _T_2197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4018;
  reg [31:0] _T_2198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4019;
  reg [31:0] _T_2198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4020;
  reg [31:0] _T_2199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4021;
  reg [31:0] _T_2199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4022;
  reg [31:0] _T_2200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4023;
  reg [31:0] _T_2200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4024;
  reg [31:0] _T_2201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4025;
  reg [31:0] _T_2201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4026;
  reg [31:0] _T_2202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4027;
  reg [31:0] _T_2202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4028;
  reg [31:0] _T_2203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4029;
  reg [31:0] _T_2203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4030;
  reg [31:0] _T_2204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4031;
  reg [31:0] _T_2204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4032;
  reg [31:0] _T_2205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4033;
  reg [31:0] _T_2205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4034;
  reg [31:0] _T_2206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4035;
  reg [31:0] _T_2206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4036;
  reg [31:0] _T_2207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4037;
  reg [31:0] _T_2207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4038;
  reg [31:0] _T_2208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4039;
  reg [31:0] _T_2208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4040;
  reg [31:0] _T_2209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4041;
  reg [31:0] _T_2209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4042;
  reg [31:0] _T_2210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4043;
  reg [31:0] _T_2210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4044;
  reg [31:0] _T_2211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4045;
  reg [31:0] _T_2211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4046;
  reg [31:0] _T_2212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4047;
  reg [31:0] _T_2212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4048;
  reg [31:0] _T_2213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4049;
  reg [31:0] _T_2213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4050;
  reg [31:0] _T_2214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4051;
  reg [31:0] _T_2214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4052;
  reg [31:0] _T_2215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4053;
  reg [31:0] _T_2215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4054;
  reg [31:0] _T_2216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4055;
  reg [31:0] _T_2216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4056;
  reg [31:0] _T_2217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4057;
  reg [31:0] _T_2217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4058;
  reg [31:0] _T_2218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4059;
  reg [31:0] _T_2218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4060;
  reg [31:0] _T_2219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4061;
  reg [31:0] _T_2219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4062;
  reg [31:0] _T_2220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4063;
  reg [31:0] _T_2220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4064;
  reg [31:0] _T_2221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4065;
  reg [31:0] _T_2221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4066;
  reg [31:0] _T_2222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4067;
  reg [31:0] _T_2222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4068;
  reg [31:0] _T_2223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4069;
  reg [31:0] _T_2223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4070;
  reg [31:0] _T_2224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4071;
  reg [31:0] _T_2224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4072;
  reg [31:0] _T_2225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4073;
  reg [31:0] _T_2225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4074;
  reg [31:0] _T_2226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4075;
  reg [31:0] _T_2226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4076;
  reg [31:0] _T_2227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4077;
  reg [31:0] _T_2227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4078;
  reg [31:0] _T_2228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4079;
  reg [31:0] _T_2228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4080;
  reg [31:0] _T_2229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4081;
  reg [31:0] _T_2229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4082;
  reg [31:0] _T_2230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4083;
  reg [31:0] _T_2230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4084;
  reg [31:0] _T_2231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4085;
  reg [31:0] _T_2231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4086;
  reg [31:0] _T_2232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4087;
  reg [31:0] _T_2232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4088;
  reg [31:0] _T_2233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4089;
  reg [31:0] _T_2233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4090;
  reg [31:0] _T_2234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4091;
  reg [31:0] _T_2234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4092;
  reg [31:0] _T_2235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4093;
  reg [31:0] _T_2235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4094;
  reg [31:0] _T_2236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4095;
  reg [31:0] _T_2236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4096;
  reg [31:0] _T_2237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4097;
  reg [31:0] _T_2237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4098;
  reg [31:0] _T_2238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4099;
  reg [31:0] _T_2238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4100;
  reg [31:0] _T_2239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4101;
  reg [31:0] _T_2239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4102;
  reg [31:0] _T_2242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4103;
  reg [31:0] _T_2242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4104;
  reg [31:0] _T_2243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4105;
  reg [31:0] _T_2243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4106;
  reg [31:0] _T_2244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4107;
  reg [31:0] _T_2244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4108;
  reg [31:0] _T_2245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4109;
  reg [31:0] _T_2245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4110;
  reg [31:0] _T_2246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4111;
  reg [31:0] _T_2246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4112;
  reg [31:0] _T_2247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4113;
  reg [31:0] _T_2247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4114;
  reg [31:0] _T_2248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4115;
  reg [31:0] _T_2248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4116;
  reg [31:0] _T_2249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4117;
  reg [31:0] _T_2249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4118;
  reg [31:0] _T_2250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4119;
  reg [31:0] _T_2250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4120;
  reg [31:0] _T_2251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4121;
  reg [31:0] _T_2251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4122;
  reg [31:0] _T_2252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4123;
  reg [31:0] _T_2252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4124;
  reg [31:0] _T_2253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4125;
  reg [31:0] _T_2253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4126;
  reg [31:0] _T_2254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4127;
  reg [31:0] _T_2254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4128;
  reg [31:0] _T_2255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4129;
  reg [31:0] _T_2255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4130;
  reg [31:0] _T_2256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4131;
  reg [31:0] _T_2256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4132;
  reg [31:0] _T_2257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4133;
  reg [31:0] _T_2257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4134;
  reg [31:0] _T_2258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4135;
  reg [31:0] _T_2258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4136;
  reg [31:0] _T_2259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4137;
  reg [31:0] _T_2259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4138;
  reg [31:0] _T_2260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4139;
  reg [31:0] _T_2260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4140;
  reg [31:0] _T_2261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4141;
  reg [31:0] _T_2261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4142;
  reg [31:0] _T_2262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4143;
  reg [31:0] _T_2262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4144;
  reg [31:0] _T_2263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4145;
  reg [31:0] _T_2263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4146;
  reg [31:0] _T_2264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4147;
  reg [31:0] _T_2264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4148;
  reg [31:0] _T_2265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4149;
  reg [31:0] _T_2265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4150;
  reg [31:0] _T_2266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4151;
  reg [31:0] _T_2266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4152;
  reg [31:0] _T_2267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4153;
  reg [31:0] _T_2267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4154;
  reg [31:0] _T_2268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4155;
  reg [31:0] _T_2268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4156;
  reg [31:0] _T_2269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4157;
  reg [31:0] _T_2269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4158;
  reg [31:0] _T_2270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4159;
  reg [31:0] _T_2270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4160;
  reg [31:0] _T_2271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4161;
  reg [31:0] _T_2271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4162;
  reg [31:0] _T_2272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4163;
  reg [31:0] _T_2272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4164;
  reg [31:0] _T_2273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4165;
  reg [31:0] _T_2273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4166;
  reg [31:0] _T_2274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4167;
  reg [31:0] _T_2274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4168;
  reg [31:0] _T_2275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4169;
  reg [31:0] _T_2275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4170;
  reg [31:0] _T_2276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4171;
  reg [31:0] _T_2276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4172;
  reg [31:0] _T_2277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4173;
  reg [31:0] _T_2277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4174;
  reg [31:0] _T_2278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4175;
  reg [31:0] _T_2278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4176;
  reg [31:0] _T_2279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4177;
  reg [31:0] _T_2279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4178;
  reg [31:0] _T_2280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4179;
  reg [31:0] _T_2280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4180;
  reg [31:0] _T_2281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4181;
  reg [31:0] _T_2281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4182;
  reg [31:0] _T_2282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4183;
  reg [31:0] _T_2282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4184;
  reg [31:0] _T_2283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4185;
  reg [31:0] _T_2283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4186;
  reg [31:0] _T_2284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4187;
  reg [31:0] _T_2284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4188;
  reg [31:0] _T_2285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4189;
  reg [31:0] _T_2285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4190;
  reg [31:0] _T_2286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4191;
  reg [31:0] _T_2286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4192;
  reg [31:0] _T_2287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4193;
  reg [31:0] _T_2287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4194;
  reg [31:0] _T_2288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4195;
  reg [31:0] _T_2288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4196;
  reg [31:0] _T_2289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4197;
  reg [31:0] _T_2289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4198;
  reg [31:0] _T_2290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4199;
  reg [31:0] _T_2290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4200;
  reg [31:0] _T_2291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4201;
  reg [31:0] _T_2291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4202;
  reg [31:0] _T_2292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4203;
  reg [31:0] _T_2292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4204;
  reg [31:0] _T_2293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4205;
  reg [31:0] _T_2293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4206;
  reg [31:0] _T_2294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4207;
  reg [31:0] _T_2294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4208;
  reg [31:0] _T_2295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4209;
  reg [31:0] _T_2295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4210;
  reg [31:0] _T_2296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4211;
  reg [31:0] _T_2296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4212;
  reg [31:0] _T_2297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4213;
  reg [31:0] _T_2297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4214;
  reg [31:0] _T_2298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4215;
  reg [31:0] _T_2298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4216;
  reg [31:0] _T_2299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4217;
  reg [31:0] _T_2299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4218;
  reg [31:0] _T_2300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4219;
  reg [31:0] _T_2300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4220;
  reg [31:0] _T_2301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4221;
  reg [31:0] _T_2301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4222;
  reg [31:0] _T_2302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4223;
  reg [31:0] _T_2302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4224;
  reg [31:0] _T_2303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4225;
  reg [31:0] _T_2303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4226;
  reg [31:0] _T_2304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4227;
  reg [31:0] _T_2304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4228;
  reg [31:0] _T_2305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4229;
  reg [31:0] _T_2305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4230;
  reg [31:0] _T_2306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4231;
  reg [31:0] _T_2306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4232;
  reg [31:0] _T_2307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4233;
  reg [31:0] _T_2307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4234;
  reg [31:0] _T_2308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4235;
  reg [31:0] _T_2308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4236;
  reg [31:0] _T_2309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4237;
  reg [31:0] _T_2309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4238;
  reg [31:0] _T_2310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4239;
  reg [31:0] _T_2310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4240;
  reg [31:0] _T_2311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4241;
  reg [31:0] _T_2311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4242;
  reg [31:0] _T_2312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4243;
  reg [31:0] _T_2312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4244;
  reg [31:0] _T_2313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4245;
  reg [31:0] _T_2313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4246;
  reg [31:0] _T_2314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4247;
  reg [31:0] _T_2314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4248;
  reg [31:0] _T_2315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4249;
  reg [31:0] _T_2315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4250;
  reg [31:0] _T_2316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4251;
  reg [31:0] _T_2316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4252;
  reg [31:0] _T_2317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4253;
  reg [31:0] _T_2317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4254;
  reg [31:0] _T_2318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4255;
  reg [31:0] _T_2318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4256;
  reg [31:0] _T_2319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4257;
  reg [31:0] _T_2319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4258;
  reg [31:0] _T_2320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4259;
  reg [31:0] _T_2320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4260;
  reg [31:0] _T_2321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4261;
  reg [31:0] _T_2321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4262;
  reg [31:0] _T_2322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4263;
  reg [31:0] _T_2322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4264;
  reg [31:0] _T_2323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4265;
  reg [31:0] _T_2323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4266;
  reg [31:0] _T_2324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4267;
  reg [31:0] _T_2324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4268;
  reg [31:0] _T_2325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4269;
  reg [31:0] _T_2325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4270;
  reg [31:0] _T_2326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4271;
  reg [31:0] _T_2326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4272;
  reg [31:0] _T_2327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4273;
  reg [31:0] _T_2327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4274;
  reg [31:0] _T_2328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4275;
  reg [31:0] _T_2328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4276;
  reg [31:0] _T_2329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4277;
  reg [31:0] _T_2329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4278;
  reg [31:0] _T_2330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4279;
  reg [31:0] _T_2330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4280;
  reg [31:0] _T_2331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4281;
  reg [31:0] _T_2331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4282;
  reg [31:0] _T_2332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4283;
  reg [31:0] _T_2332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4284;
  reg [31:0] _T_2333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4285;
  reg [31:0] _T_2333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4286;
  reg [31:0] _T_2334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4287;
  reg [31:0] _T_2334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4288;
  reg [31:0] _T_2335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4289;
  reg [31:0] _T_2335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4290;
  reg [31:0] _T_2336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4291;
  reg [31:0] _T_2336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4292;
  reg [31:0] _T_2337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4293;
  reg [31:0] _T_2337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4294;
  reg [31:0] _T_2338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4295;
  reg [31:0] _T_2338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4296;
  reg [31:0] _T_2339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4297;
  reg [31:0] _T_2339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4298;
  reg [31:0] _T_2340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4299;
  reg [31:0] _T_2340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4300;
  reg [31:0] _T_2341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4301;
  reg [31:0] _T_2341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4302;
  reg [31:0] _T_2342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4303;
  reg [31:0] _T_2342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4304;
  reg [31:0] _T_2343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4305;
  reg [31:0] _T_2343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4306;
  reg [31:0] _T_2344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4307;
  reg [31:0] _T_2344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4308;
  reg [31:0] _T_2345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4309;
  reg [31:0] _T_2345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4310;
  reg [31:0] _T_2346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4311;
  reg [31:0] _T_2346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4312;
  reg [31:0] _T_2347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4313;
  reg [31:0] _T_2347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4314;
  reg [31:0] _T_2348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4315;
  reg [31:0] _T_2348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4316;
  reg [31:0] _T_2349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4317;
  reg [31:0] _T_2349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4318;
  reg [31:0] _T_2350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4319;
  reg [31:0] _T_2350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4320;
  reg [31:0] _T_2351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4321;
  reg [31:0] _T_2351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4322;
  reg [31:0] _T_2352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4323;
  reg [31:0] _T_2352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4324;
  reg [31:0] _T_2353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4325;
  reg [31:0] _T_2353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4326;
  reg [31:0] _T_2354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4327;
  reg [31:0] _T_2354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4328;
  reg [31:0] _T_2355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4329;
  reg [31:0] _T_2355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4330;
  reg [31:0] _T_2356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4331;
  reg [31:0] _T_2356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4332;
  reg [31:0] _T_2357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4333;
  reg [31:0] _T_2357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4334;
  reg [31:0] _T_2358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4335;
  reg [31:0] _T_2358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4336;
  reg [31:0] _T_2359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4337;
  reg [31:0] _T_2359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4338;
  reg [31:0] _T_2360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4339;
  reg [31:0] _T_2360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4340;
  reg [31:0] _T_2361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4341;
  reg [31:0] _T_2361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4342;
  reg [31:0] _T_2362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4343;
  reg [31:0] _T_2362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4344;
  reg [31:0] _T_2363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4345;
  reg [31:0] _T_2363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4346;
  reg [31:0] _T_2364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4347;
  reg [31:0] _T_2364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4348;
  reg [31:0] _T_2365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4349;
  reg [31:0] _T_2365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4350;
  reg [31:0] _T_2366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4351;
  reg [31:0] _T_2366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4352;
  reg [31:0] _T_2367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4353;
  reg [31:0] _T_2367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4354;
  reg [31:0] _T_2368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4355;
  reg [31:0] _T_2368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4356;
  reg [31:0] _T_2369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4357;
  reg [31:0] _T_2369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4358;
  reg [31:0] _T_2370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4359;
  reg [31:0] _T_2370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4360;
  reg [31:0] _T_2371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4361;
  reg [31:0] _T_2371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4362;
  reg [31:0] _T_2372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4363;
  reg [31:0] _T_2372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4364;
  reg [31:0] _T_2373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4365;
  reg [31:0] _T_2373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4366;
  reg [31:0] _T_2374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4367;
  reg [31:0] _T_2374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4368;
  reg [31:0] _T_2375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4369;
  reg [31:0] _T_2375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4370;
  reg [31:0] _T_2376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4371;
  reg [31:0] _T_2376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4372;
  reg [31:0] _T_2377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4373;
  reg [31:0] _T_2377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4374;
  reg [31:0] _T_2378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4375;
  reg [31:0] _T_2378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4376;
  reg [31:0] _T_2379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4377;
  reg [31:0] _T_2379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4378;
  reg [31:0] _T_2380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4379;
  reg [31:0] _T_2380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4380;
  reg [31:0] _T_2381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4381;
  reg [31:0] _T_2381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4382;
  reg [31:0] _T_2382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4383;
  reg [31:0] _T_2382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4384;
  reg [31:0] _T_2383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4385;
  reg [31:0] _T_2383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4386;
  reg [31:0] _T_2384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4387;
  reg [31:0] _T_2384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4388;
  reg [31:0] _T_2385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4389;
  reg [31:0] _T_2385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4390;
  reg [31:0] _T_2386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4391;
  reg [31:0] _T_2386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4392;
  reg [31:0] _T_2387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4393;
  reg [31:0] _T_2387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4394;
  reg [31:0] _T_2388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4395;
  reg [31:0] _T_2388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4396;
  reg [31:0] _T_2389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4397;
  reg [31:0] _T_2389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4398;
  reg [31:0] _T_2390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4399;
  reg [31:0] _T_2390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4400;
  reg [31:0] _T_2391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4401;
  reg [31:0] _T_2391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4402;
  reg [31:0] _T_2392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4403;
  reg [31:0] _T_2392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4404;
  reg [31:0] _T_2393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4405;
  reg [31:0] _T_2393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4406;
  reg [31:0] _T_2394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4407;
  reg [31:0] _T_2394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4408;
  reg [31:0] _T_2395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4409;
  reg [31:0] _T_2395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4410;
  reg [31:0] _T_2396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4411;
  reg [31:0] _T_2396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4412;
  reg [31:0] _T_2397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4413;
  reg [31:0] _T_2397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4414;
  reg [31:0] _T_2398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4415;
  reg [31:0] _T_2398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4416;
  reg [31:0] _T_2399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4417;
  reg [31:0] _T_2399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4418;
  reg [31:0] _T_2400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4419;
  reg [31:0] _T_2400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4420;
  reg [31:0] _T_2401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4421;
  reg [31:0] _T_2401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4422;
  reg [31:0] _T_2402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4423;
  reg [31:0] _T_2402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4424;
  reg [31:0] _T_2403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4425;
  reg [31:0] _T_2403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4426;
  reg [31:0] _T_2404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4427;
  reg [31:0] _T_2404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4428;
  reg [31:0] _T_2405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4429;
  reg [31:0] _T_2405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4430;
  reg [31:0] _T_2406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4431;
  reg [31:0] _T_2406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4432;
  reg [31:0] _T_2407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4433;
  reg [31:0] _T_2407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4434;
  reg [31:0] _T_2408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4435;
  reg [31:0] _T_2408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4436;
  reg [31:0] _T_2409_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4437;
  reg [31:0] _T_2409_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4438;
  reg [31:0] _T_2410_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4439;
  reg [31:0] _T_2410_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4440;
  reg [31:0] _T_2411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4441;
  reg [31:0] _T_2411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4442;
  reg [31:0] _T_2412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4443;
  reg [31:0] _T_2412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4444;
  reg [31:0] _T_2413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4445;
  reg [31:0] _T_2413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4446;
  reg [31:0] _T_2414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4447;
  reg [31:0] _T_2414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4448;
  reg [31:0] _T_2415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4449;
  reg [31:0] _T_2415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4450;
  reg [31:0] _T_2416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4451;
  reg [31:0] _T_2416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4452;
  reg [31:0] _T_2417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4453;
  reg [31:0] _T_2417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4454;
  reg [31:0] _T_2418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4455;
  reg [31:0] _T_2418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4456;
  reg [31:0] _T_2419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4457;
  reg [31:0] _T_2419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4458;
  reg [31:0] _T_2420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4459;
  reg [31:0] _T_2420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4460;
  reg [31:0] _T_2421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4461;
  reg [31:0] _T_2421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4462;
  reg [31:0] _T_2422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4463;
  reg [31:0] _T_2422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4464;
  reg [31:0] _T_2423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4465;
  reg [31:0] _T_2423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4466;
  reg [31:0] _T_2424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4467;
  reg [31:0] _T_2424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4468;
  reg [31:0] _T_2425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4469;
  reg [31:0] _T_2425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4470;
  reg [31:0] _T_2426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4471;
  reg [31:0] _T_2426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4472;
  reg [31:0] _T_2427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4473;
  reg [31:0] _T_2427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4474;
  reg [31:0] _T_2428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4475;
  reg [31:0] _T_2428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4476;
  reg [31:0] _T_2429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4477;
  reg [31:0] _T_2429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4478;
  reg [31:0] _T_2430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4479;
  reg [31:0] _T_2430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4480;
  reg [31:0] _T_2431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4481;
  reg [31:0] _T_2431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4482;
  reg [31:0] _T_2432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4483;
  reg [31:0] _T_2432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4484;
  reg [31:0] _T_2433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4485;
  reg [31:0] _T_2433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4486;
  reg [31:0] _T_2434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4487;
  reg [31:0] _T_2434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4488;
  reg [31:0] _T_2435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4489;
  reg [31:0] _T_2435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4490;
  reg [31:0] _T_2436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4491;
  reg [31:0] _T_2436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4492;
  reg [31:0] _T_2437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4493;
  reg [31:0] _T_2437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4494;
  reg [31:0] _T_2438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4495;
  reg [31:0] _T_2438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4496;
  reg [31:0] _T_2439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4497;
  reg [31:0] _T_2439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4498;
  reg [31:0] _T_2440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4499;
  reg [31:0] _T_2440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4500;
  reg [31:0] _T_2441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4501;
  reg [31:0] _T_2441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4502;
  reg [31:0] _T_2442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4503;
  reg [31:0] _T_2442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4504;
  reg [31:0] _T_2443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4505;
  reg [31:0] _T_2443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4506;
  reg [31:0] _T_2444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4507;
  reg [31:0] _T_2444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4508;
  reg [31:0] _T_2445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4509;
  reg [31:0] _T_2445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4510;
  reg [31:0] _T_2446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4511;
  reg [31:0] _T_2446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4512;
  reg [31:0] _T_2447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4513;
  reg [31:0] _T_2447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4514;
  reg [31:0] _T_2448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4515;
  reg [31:0] _T_2448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4516;
  reg [31:0] _T_2449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4517;
  reg [31:0] _T_2449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4518;
  reg [31:0] _T_2450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4519;
  reg [31:0] _T_2450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4520;
  reg [31:0] _T_2451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4521;
  reg [31:0] _T_2451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4522;
  reg [31:0] _T_2452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4523;
  reg [31:0] _T_2452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4524;
  reg [31:0] _T_2453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4525;
  reg [31:0] _T_2453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4526;
  reg [31:0] _T_2454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4527;
  reg [31:0] _T_2454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4528;
  reg [31:0] _T_2455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4529;
  reg [31:0] _T_2455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4530;
  reg [31:0] _T_2456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4531;
  reg [31:0] _T_2456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4532;
  reg [31:0] _T_2457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4533;
  reg [31:0] _T_2457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4534;
  reg [31:0] _T_2458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4535;
  reg [31:0] _T_2458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4536;
  reg [31:0] _T_2459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4537;
  reg [31:0] _T_2459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4538;
  reg [31:0] _T_2460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4539;
  reg [31:0] _T_2460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4540;
  reg [31:0] _T_2461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4541;
  reg [31:0] _T_2461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4542;
  reg [31:0] _T_2462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4543;
  reg [31:0] _T_2462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4544;
  reg [31:0] _T_2463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4545;
  reg [31:0] _T_2463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4546;
  reg [31:0] _T_2464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4547;
  reg [31:0] _T_2464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4548;
  reg [31:0] _T_2465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4549;
  reg [31:0] _T_2465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4550;
  reg [31:0] _T_2466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4551;
  reg [31:0] _T_2466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4552;
  reg [31:0] _T_2467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4553;
  reg [31:0] _T_2467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4554;
  reg [31:0] _T_2468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4555;
  reg [31:0] _T_2468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4556;
  reg [31:0] _T_2469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4557;
  reg [31:0] _T_2469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4558;
  reg [31:0] _T_2470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4559;
  reg [31:0] _T_2470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4560;
  reg [31:0] _T_2471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4561;
  reg [31:0] _T_2471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4562;
  reg [31:0] _T_2472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4563;
  reg [31:0] _T_2472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4564;
  reg [31:0] _T_2473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4565;
  reg [31:0] _T_2473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4566;
  reg [31:0] _T_2474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4567;
  reg [31:0] _T_2474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4568;
  reg [31:0] _T_2475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4569;
  reg [31:0] _T_2475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4570;
  reg [31:0] _T_2476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4571;
  reg [31:0] _T_2476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4572;
  reg [31:0] _T_2477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4573;
  reg [31:0] _T_2477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4574;
  reg [31:0] _T_2478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4575;
  reg [31:0] _T_2478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4576;
  reg [31:0] _T_2479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4577;
  reg [31:0] _T_2479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4578;
  reg [31:0] _T_2480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4579;
  reg [31:0] _T_2480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4580;
  reg [31:0] _T_2481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4581;
  reg [31:0] _T_2481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4582;
  reg [31:0] _T_2482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4583;
  reg [31:0] _T_2482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4584;
  reg [31:0] _T_2483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4585;
  reg [31:0] _T_2483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4586;
  reg [31:0] _T_2484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4587;
  reg [31:0] _T_2484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4588;
  reg [31:0] _T_2485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4589;
  reg [31:0] _T_2485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4590;
  reg [31:0] _T_2486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4591;
  reg [31:0] _T_2486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4592;
  reg [31:0] _T_2487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4593;
  reg [31:0] _T_2487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4594;
  reg [31:0] _T_2488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4595;
  reg [31:0] _T_2488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4596;
  reg [31:0] _T_2489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4597;
  reg [31:0] _T_2489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4598;
  reg [31:0] _T_2490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4599;
  reg [31:0] _T_2490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4600;
  reg [31:0] _T_2491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4601;
  reg [31:0] _T_2491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4602;
  reg [31:0] _T_2492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4603;
  reg [31:0] _T_2492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4604;
  reg [31:0] _T_2493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4605;
  reg [31:0] _T_2493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4606;
  reg [31:0] _T_2494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4607;
  reg [31:0] _T_2494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4608;
  reg [31:0] _T_2495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4609;
  reg [31:0] _T_2495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4610;
  reg [31:0] _T_2496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4611;
  reg [31:0] _T_2496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4612;
  reg [31:0] _T_2497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4613;
  reg [31:0] _T_2497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4614;
  wire [63:0] _T_2502;
  reg [31:0] _T_2507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4615;
  reg [31:0] _T_2507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4616;
  reg [31:0] _T_2508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4617;
  reg [31:0] _T_2508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4618;
  reg [31:0] _T_2509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4619;
  reg [31:0] _T_2509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4620;
  reg [31:0] _T_2510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4621;
  reg [31:0] _T_2510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4622;
  reg [31:0] _T_2511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4623;
  reg [31:0] _T_2511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4624;
  reg [31:0] _T_2512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4625;
  reg [31:0] _T_2512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4626;
  reg [31:0] _T_2513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4627;
  reg [31:0] _T_2513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4628;
  reg [31:0] _T_2514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4629;
  reg [31:0] _T_2514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4630;
  reg [31:0] _T_2515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4631;
  reg [31:0] _T_2515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4632;
  reg [31:0] _T_2516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4633;
  reg [31:0] _T_2516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4634;
  reg [31:0] _T_2517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4635;
  reg [31:0] _T_2517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4636;
  reg [31:0] _T_2518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4637;
  reg [31:0] _T_2518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4638;
  reg [31:0] _T_2519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4639;
  reg [31:0] _T_2519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4640;
  reg [31:0] _T_2520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4641;
  reg [31:0] _T_2520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4642;
  reg [31:0] _T_2521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4643;
  reg [31:0] _T_2521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4644;
  reg [31:0] _T_2522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4645;
  reg [31:0] _T_2522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4646;
  reg [31:0] _T_2523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4647;
  reg [31:0] _T_2523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4648;
  reg [31:0] _T_2524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4649;
  reg [31:0] _T_2524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4650;
  reg [31:0] _T_2525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4651;
  reg [31:0] _T_2525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4652;
  reg [31:0] _T_2526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4653;
  reg [31:0] _T_2526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4654;
  reg [31:0] _T_2527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4655;
  reg [31:0] _T_2527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4656;
  reg [31:0] _T_2528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4657;
  reg [31:0] _T_2528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4658;
  reg [31:0] _T_2529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4659;
  reg [31:0] _T_2529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4660;
  reg [31:0] _T_2530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4661;
  reg [31:0] _T_2530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4662;
  reg [31:0] _T_2531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4663;
  reg [31:0] _T_2531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4664;
  reg [31:0] _T_2532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4665;
  reg [31:0] _T_2532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4666;
  reg [31:0] _T_2533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4667;
  reg [31:0] _T_2533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4668;
  reg [31:0] _T_2534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4669;
  reg [31:0] _T_2534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4670;
  reg [31:0] _T_2535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4671;
  reg [31:0] _T_2535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4672;
  reg [31:0] _T_2536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4673;
  reg [31:0] _T_2536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4674;
  reg [31:0] _T_2537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4675;
  reg [31:0] _T_2537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4676;
  reg [31:0] _T_2538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4677;
  reg [31:0] _T_2538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4678;
  reg [31:0] _T_2539_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4679;
  reg [31:0] _T_2539_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4680;
  reg [31:0] _T_2540_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4681;
  reg [31:0] _T_2540_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4682;
  reg [31:0] _T_2541_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4683;
  reg [31:0] _T_2541_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4684;
  reg [31:0] _T_2542_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4685;
  reg [31:0] _T_2542_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4686;
  reg [31:0] _T_2543_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4687;
  reg [31:0] _T_2543_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4688;
  reg [31:0] _T_2544_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4689;
  reg [31:0] _T_2544_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4690;
  reg [31:0] _T_2545_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4691;
  reg [31:0] _T_2545_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4692;
  reg [31:0] _T_2546_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4693;
  reg [31:0] _T_2546_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4694;
  reg [31:0] _T_2547_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4695;
  reg [31:0] _T_2547_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4696;
  reg [31:0] _T_2548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4697;
  reg [31:0] _T_2548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4698;
  reg [31:0] _T_2549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4699;
  reg [31:0] _T_2549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4700;
  reg [31:0] _T_2550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4701;
  reg [31:0] _T_2550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4702;
  reg [31:0] _T_2551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4703;
  reg [31:0] _T_2551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4704;
  reg [31:0] _T_2552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4705;
  reg [31:0] _T_2552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4706;
  reg [31:0] _T_2553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4707;
  reg [31:0] _T_2553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4708;
  reg [31:0] _T_2554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4709;
  reg [31:0] _T_2554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4710;
  reg [31:0] _T_2555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4711;
  reg [31:0] _T_2555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4712;
  reg [31:0] _T_2556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4713;
  reg [31:0] _T_2556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4714;
  reg [31:0] _T_2557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4715;
  reg [31:0] _T_2557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4716;
  reg [31:0] _T_2558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4717;
  reg [31:0] _T_2558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4718;
  reg [31:0] _T_2559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4719;
  reg [31:0] _T_2559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4720;
  reg [31:0] _T_2560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4721;
  reg [31:0] _T_2560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4722;
  reg [31:0] _T_2561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4723;
  reg [31:0] _T_2561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4724;
  reg [31:0] _T_2562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4725;
  reg [31:0] _T_2562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4726;
  reg [31:0] _T_2563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4727;
  reg [31:0] _T_2563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4728;
  reg [31:0] _T_2564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4729;
  reg [31:0] _T_2564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4730;
  reg [31:0] _T_2565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4731;
  reg [31:0] _T_2565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4732;
  reg [31:0] _T_2566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4733;
  reg [31:0] _T_2566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4734;
  reg [31:0] _T_2567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4735;
  reg [31:0] _T_2567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4736;
  reg [31:0] _T_2568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4737;
  reg [31:0] _T_2568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4738;
  reg [31:0] _T_2569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4739;
  reg [31:0] _T_2569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4740;
  reg [31:0] _T_2570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4741;
  reg [31:0] _T_2570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4742;
  reg [31:0] _T_2571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4743;
  reg [31:0] _T_2571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4744;
  reg [31:0] _T_2572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4745;
  reg [31:0] _T_2572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4746;
  reg [31:0] _T_2573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4747;
  reg [31:0] _T_2573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4748;
  reg [31:0] _T_2574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4749;
  reg [31:0] _T_2574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4750;
  reg [31:0] _T_2575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4751;
  reg [31:0] _T_2575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4752;
  reg [31:0] _T_2576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4753;
  reg [31:0] _T_2576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4754;
  reg [31:0] _T_2577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4755;
  reg [31:0] _T_2577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4756;
  reg [31:0] _T_2578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4757;
  reg [31:0] _T_2578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4758;
  reg [31:0] _T_2579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4759;
  reg [31:0] _T_2579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4760;
  reg [31:0] _T_2580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4761;
  reg [31:0] _T_2580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4762;
  reg [31:0] _T_2581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4763;
  reg [31:0] _T_2581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4764;
  reg [31:0] _T_2582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4765;
  reg [31:0] _T_2582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4766;
  reg [31:0] _T_2583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4767;
  reg [31:0] _T_2583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4768;
  reg [31:0] _T_2584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4769;
  reg [31:0] _T_2584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4770;
  reg [31:0] _T_2585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4771;
  reg [31:0] _T_2585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4772;
  reg [31:0] _T_2586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4773;
  reg [31:0] _T_2586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4774;
  reg [31:0] _T_2587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4775;
  reg [31:0] _T_2587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4776;
  reg [31:0] _T_2588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4777;
  reg [31:0] _T_2588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4778;
  reg [31:0] _T_2589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4779;
  reg [31:0] _T_2589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4780;
  reg [31:0] _T_2590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4781;
  reg [31:0] _T_2590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4782;
  reg [31:0] _T_2591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4783;
  reg [31:0] _T_2591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4784;
  reg [31:0] _T_2592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4785;
  reg [31:0] _T_2592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4786;
  reg [31:0] _T_2593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4787;
  reg [31:0] _T_2593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4788;
  reg [31:0] _T_2594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4789;
  reg [31:0] _T_2594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4790;
  reg [31:0] _T_2595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4791;
  reg [31:0] _T_2595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4792;
  reg [31:0] _T_2596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4793;
  reg [31:0] _T_2596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4794;
  reg [31:0] _T_2597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4795;
  reg [31:0] _T_2597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4796;
  reg [31:0] _T_2598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4797;
  reg [31:0] _T_2598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4798;
  reg [31:0] _T_2599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4799;
  reg [31:0] _T_2599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4800;
  reg [31:0] _T_2600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4801;
  reg [31:0] _T_2600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4802;
  reg [31:0] _T_2601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4803;
  reg [31:0] _T_2601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4804;
  reg [31:0] _T_2602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4805;
  reg [31:0] _T_2602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4806;
  reg [31:0] _T_2603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4807;
  reg [31:0] _T_2603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4808;
  reg [31:0] _T_2604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4809;
  reg [31:0] _T_2604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4810;
  reg [31:0] _T_2605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4811;
  reg [31:0] _T_2605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4812;
  reg [31:0] _T_2606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4813;
  reg [31:0] _T_2606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4814;
  reg [31:0] _T_2607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4815;
  reg [31:0] _T_2607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4816;
  reg [31:0] _T_2608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4817;
  reg [31:0] _T_2608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4818;
  reg [31:0] _T_2609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4819;
  reg [31:0] _T_2609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4820;
  reg [31:0] _T_2610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4821;
  reg [31:0] _T_2610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4822;
  reg [31:0] _T_2611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4823;
  reg [31:0] _T_2611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4824;
  reg [31:0] _T_2612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4825;
  reg [31:0] _T_2612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4826;
  reg [31:0] _T_2613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4827;
  reg [31:0] _T_2613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4828;
  reg [31:0] _T_2614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4829;
  reg [31:0] _T_2614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4830;
  reg [31:0] _T_2615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4831;
  reg [31:0] _T_2615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4832;
  reg [31:0] _T_2616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4833;
  reg [31:0] _T_2616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4834;
  reg [31:0] _T_2617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4835;
  reg [31:0] _T_2617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4836;
  reg [31:0] _T_2618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4837;
  reg [31:0] _T_2618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4838;
  reg [31:0] _T_2619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4839;
  reg [31:0] _T_2619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4840;
  reg [31:0] _T_2620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4841;
  reg [31:0] _T_2620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4842;
  reg [31:0] _T_2621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4843;
  reg [31:0] _T_2621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4844;
  reg [31:0] _T_2622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4845;
  reg [31:0] _T_2622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4846;
  reg [31:0] _T_2623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4847;
  reg [31:0] _T_2623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4848;
  reg [31:0] _T_2624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4849;
  reg [31:0] _T_2624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4850;
  reg [31:0] _T_2625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4851;
  reg [31:0] _T_2625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4852;
  reg [31:0] _T_2626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4853;
  reg [31:0] _T_2626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4854;
  reg [31:0] _T_2627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4855;
  reg [31:0] _T_2627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4856;
  reg [31:0] _T_2628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4857;
  reg [31:0] _T_2628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4858;
  reg [31:0] _T_2629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4859;
  reg [31:0] _T_2629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4860;
  reg [31:0] _T_2630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4861;
  reg [31:0] _T_2630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4862;
  reg [31:0] _T_2631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4863;
  reg [31:0] _T_2631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4864;
  reg [31:0] _T_2632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4865;
  reg [31:0] _T_2632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4866;
  reg [31:0] _T_2633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4867;
  reg [31:0] _T_2633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4868;
  reg [31:0] _T_2634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4869;
  reg [31:0] _T_2634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4870;
  reg [31:0] _T_2635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4871;
  reg [31:0] _T_2635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4872;
  reg [31:0] _T_2636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4873;
  reg [31:0] _T_2636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4874;
  reg [31:0] _T_2637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4875;
  reg [31:0] _T_2637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4876;
  reg [31:0] _T_2638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4877;
  reg [31:0] _T_2638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4878;
  reg [31:0] _T_2639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4879;
  reg [31:0] _T_2639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4880;
  reg [31:0] _T_2640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4881;
  reg [31:0] _T_2640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4882;
  reg [31:0] _T_2641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4883;
  reg [31:0] _T_2641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4884;
  reg [31:0] _T_2642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4885;
  reg [31:0] _T_2642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4886;
  reg [31:0] _T_2643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4887;
  reg [31:0] _T_2643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4888;
  reg [31:0] _T_2644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4889;
  reg [31:0] _T_2644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4890;
  reg [31:0] _T_2645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4891;
  reg [31:0] _T_2645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4892;
  reg [31:0] _T_2646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4893;
  reg [31:0] _T_2646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4894;
  reg [31:0] _T_2647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4895;
  reg [31:0] _T_2647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4896;
  reg [31:0] _T_2648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4897;
  reg [31:0] _T_2648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4898;
  reg [31:0] _T_2649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4899;
  reg [31:0] _T_2649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4900;
  reg [31:0] _T_2650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4901;
  reg [31:0] _T_2650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4902;
  reg [31:0] _T_2651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4903;
  reg [31:0] _T_2651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4904;
  reg [31:0] _T_2652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4905;
  reg [31:0] _T_2652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4906;
  reg [31:0] _T_2653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4907;
  reg [31:0] _T_2653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4908;
  reg [31:0] _T_2654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4909;
  reg [31:0] _T_2654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4910;
  reg [31:0] _T_2655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4911;
  reg [31:0] _T_2655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4912;
  reg [31:0] _T_2656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4913;
  reg [31:0] _T_2656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4914;
  reg [31:0] _T_2657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4915;
  reg [31:0] _T_2657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4916;
  reg [31:0] _T_2658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4917;
  reg [31:0] _T_2658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4918;
  reg [31:0] _T_2659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4919;
  reg [31:0] _T_2659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4920;
  reg [31:0] _T_2660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4921;
  reg [31:0] _T_2660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4922;
  reg [31:0] _T_2661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4923;
  reg [31:0] _T_2661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4924;
  reg [31:0] _T_2662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4925;
  reg [31:0] _T_2662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4926;
  reg [31:0] _T_2663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4927;
  reg [31:0] _T_2663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4928;
  reg [31:0] _T_2664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4929;
  reg [31:0] _T_2664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4930;
  reg [31:0] _T_2665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4931;
  reg [31:0] _T_2665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4932;
  reg [31:0] _T_2666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4933;
  reg [31:0] _T_2666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4934;
  reg [31:0] _T_2667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4935;
  reg [31:0] _T_2667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4936;
  reg [31:0] _T_2668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4937;
  reg [31:0] _T_2668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4938;
  reg [31:0] _T_2669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4939;
  reg [31:0] _T_2669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4940;
  reg [31:0] _T_2670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4941;
  reg [31:0] _T_2670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4942;
  reg [31:0] _T_2671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4943;
  reg [31:0] _T_2671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4944;
  reg [31:0] _T_2672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4945;
  reg [31:0] _T_2672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4946;
  reg [31:0] _T_2673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4947;
  reg [31:0] _T_2673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4948;
  reg [31:0] _T_2674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4949;
  reg [31:0] _T_2674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4950;
  reg [31:0] _T_2675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4951;
  reg [31:0] _T_2675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4952;
  reg [31:0] _T_2676_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4953;
  reg [31:0] _T_2676_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4954;
  reg [31:0] _T_2677_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4955;
  reg [31:0] _T_2677_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4956;
  reg [31:0] _T_2678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4957;
  reg [31:0] _T_2678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4958;
  reg [31:0] _T_2679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4959;
  reg [31:0] _T_2679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4960;
  reg [31:0] _T_2680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4961;
  reg [31:0] _T_2680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4962;
  reg [31:0] _T_2681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4963;
  reg [31:0] _T_2681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4964;
  reg [31:0] _T_2682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4965;
  reg [31:0] _T_2682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4966;
  reg [31:0] _T_2683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4967;
  reg [31:0] _T_2683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4968;
  reg [31:0] _T_2684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4969;
  reg [31:0] _T_2684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4970;
  reg [31:0] _T_2685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4971;
  reg [31:0] _T_2685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4972;
  reg [31:0] _T_2686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4973;
  reg [31:0] _T_2686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4974;
  reg [31:0] _T_2687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4975;
  reg [31:0] _T_2687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4976;
  reg [31:0] _T_2688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4977;
  reg [31:0] _T_2688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4978;
  reg [31:0] _T_2689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4979;
  reg [31:0] _T_2689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4980;
  reg [31:0] _T_2690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4981;
  reg [31:0] _T_2690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4982;
  reg [31:0] _T_2691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4983;
  reg [31:0] _T_2691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4984;
  reg [31:0] _T_2692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4985;
  reg [31:0] _T_2692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4986;
  reg [31:0] _T_2693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4987;
  reg [31:0] _T_2693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4988;
  reg [31:0] _T_2694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4989;
  reg [31:0] _T_2694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4990;
  reg [31:0] _T_2695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4991;
  reg [31:0] _T_2695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4992;
  reg [31:0] _T_2696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4993;
  reg [31:0] _T_2696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4994;
  reg [31:0] _T_2697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4995;
  reg [31:0] _T_2697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4996;
  reg [31:0] _T_2698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4997;
  reg [31:0] _T_2698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4998;
  reg [31:0] _T_2699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4999;
  reg [31:0] _T_2699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5000;
  reg [31:0] _T_2700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5001;
  reg [31:0] _T_2700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5002;
  reg [31:0] _T_2701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5003;
  reg [31:0] _T_2701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5004;
  reg [31:0] _T_2702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5005;
  reg [31:0] _T_2702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5006;
  reg [31:0] _T_2703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5007;
  reg [31:0] _T_2703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5008;
  reg [31:0] _T_2704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5009;
  reg [31:0] _T_2704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5010;
  reg [31:0] _T_2705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5011;
  reg [31:0] _T_2705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5012;
  reg [31:0] _T_2706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5013;
  reg [31:0] _T_2706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5014;
  reg [31:0] _T_2707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5015;
  reg [31:0] _T_2707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5016;
  reg [31:0] _T_2708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5017;
  reg [31:0] _T_2708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5018;
  reg [31:0] _T_2709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5019;
  reg [31:0] _T_2709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5020;
  reg [31:0] _T_2710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5021;
  reg [31:0] _T_2710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5022;
  reg [31:0] _T_2711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5023;
  reg [31:0] _T_2711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5024;
  reg [31:0] _T_2712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5025;
  reg [31:0] _T_2712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5026;
  reg [31:0] _T_2713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5027;
  reg [31:0] _T_2713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5028;
  reg [31:0] _T_2714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5029;
  reg [31:0] _T_2714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5030;
  reg [31:0] _T_2715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5031;
  reg [31:0] _T_2715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5032;
  reg [31:0] _T_2716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5033;
  reg [31:0] _T_2716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5034;
  reg [31:0] _T_2717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5035;
  reg [31:0] _T_2717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5036;
  reg [31:0] _T_2718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5037;
  reg [31:0] _T_2718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5038;
  reg [31:0] _T_2719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5039;
  reg [31:0] _T_2719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5040;
  reg [31:0] _T_2720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5041;
  reg [31:0] _T_2720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5042;
  reg [31:0] _T_2721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5043;
  reg [31:0] _T_2721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5044;
  reg [31:0] _T_2722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5045;
  reg [31:0] _T_2722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5046;
  reg [31:0] _T_2723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5047;
  reg [31:0] _T_2723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5048;
  reg [31:0] _T_2724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5049;
  reg [31:0] _T_2724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5050;
  reg [31:0] _T_2725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5051;
  reg [31:0] _T_2725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5052;
  reg [31:0] _T_2726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5053;
  reg [31:0] _T_2726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5054;
  reg [31:0] _T_2727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5055;
  reg [31:0] _T_2727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5056;
  reg [31:0] _T_2728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5057;
  reg [31:0] _T_2728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5058;
  reg [31:0] _T_2729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5059;
  reg [31:0] _T_2729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5060;
  reg [31:0] _T_2730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5061;
  reg [31:0] _T_2730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5062;
  reg [31:0] _T_2731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5063;
  reg [31:0] _T_2731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5064;
  reg [31:0] _T_2732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5065;
  reg [31:0] _T_2732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5066;
  reg [31:0] _T_2733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5067;
  reg [31:0] _T_2733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5068;
  reg [31:0] _T_2734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5069;
  reg [31:0] _T_2734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5070;
  reg [31:0] _T_2735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5071;
  reg [31:0] _T_2735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5072;
  reg [31:0] _T_2736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5073;
  reg [31:0] _T_2736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5074;
  reg [31:0] _T_2737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5075;
  reg [31:0] _T_2737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5076;
  reg [31:0] _T_2738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5077;
  reg [31:0] _T_2738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5078;
  reg [31:0] _T_2739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5079;
  reg [31:0] _T_2739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5080;
  reg [31:0] _T_2740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5081;
  reg [31:0] _T_2740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5082;
  reg [31:0] _T_2741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5083;
  reg [31:0] _T_2741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5084;
  reg [31:0] _T_2742_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5085;
  reg [31:0] _T_2742_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5086;
  reg [31:0] _T_2743_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5087;
  reg [31:0] _T_2743_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5088;
  reg [31:0] _T_2744_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5089;
  reg [31:0] _T_2744_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5090;
  reg [31:0] _T_2745_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5091;
  reg [31:0] _T_2745_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5092;
  reg [31:0] _T_2746_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5093;
  reg [31:0] _T_2746_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5094;
  reg [31:0] _T_2747_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5095;
  reg [31:0] _T_2747_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5096;
  reg [31:0] _T_2748_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5097;
  reg [31:0] _T_2748_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5098;
  reg [31:0] _T_2749_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5099;
  reg [31:0] _T_2749_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5100;
  reg [31:0] _T_2750_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5101;
  reg [31:0] _T_2750_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5102;
  reg [31:0] _T_2751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5103;
  reg [31:0] _T_2751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5104;
  reg [31:0] _T_2752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5105;
  reg [31:0] _T_2752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5106;
  reg [31:0] _T_2753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5107;
  reg [31:0] _T_2753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5108;
  reg [31:0] _T_2754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5109;
  reg [31:0] _T_2754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5110;
  reg [31:0] _T_2755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5111;
  reg [31:0] _T_2755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5112;
  reg [31:0] _T_2756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5113;
  reg [31:0] _T_2756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5114;
  reg [31:0] _T_2757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5115;
  reg [31:0] _T_2757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5116;
  reg [31:0] _T_2758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5117;
  reg [31:0] _T_2758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5118;
  reg [31:0] _T_2759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5119;
  reg [31:0] _T_2759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5120;
  reg [31:0] _T_2760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5121;
  reg [31:0] _T_2760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5122;
  reg [31:0] _T_2761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5123;
  reg [31:0] _T_2761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5124;
  reg [31:0] _T_2762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5125;
  reg [31:0] _T_2762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5126;
  reg [31:0] _T_2765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5127;
  reg [31:0] _T_2765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5128;
  reg [31:0] _T_2766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5129;
  reg [31:0] _T_2766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5130;
  reg [31:0] _T_2767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5131;
  reg [31:0] _T_2767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5132;
  reg [31:0] _T_2768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5133;
  reg [31:0] _T_2768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5134;
  reg [31:0] _T_2769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5135;
  reg [31:0] _T_2769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5136;
  reg [31:0] _T_2770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5137;
  reg [31:0] _T_2770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5138;
  reg [31:0] _T_2771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5139;
  reg [31:0] _T_2771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5140;
  reg [31:0] _T_2772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5141;
  reg [31:0] _T_2772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5142;
  reg [31:0] _T_2773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5143;
  reg [31:0] _T_2773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5144;
  reg [31:0] _T_2774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5145;
  reg [31:0] _T_2774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5146;
  reg [31:0] _T_2775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5147;
  reg [31:0] _T_2775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5148;
  reg [31:0] _T_2776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5149;
  reg [31:0] _T_2776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5150;
  reg [31:0] _T_2777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5151;
  reg [31:0] _T_2777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5152;
  reg [31:0] _T_2778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5153;
  reg [31:0] _T_2778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5154;
  reg [31:0] _T_2779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5155;
  reg [31:0] _T_2779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5156;
  reg [31:0] _T_2780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5157;
  reg [31:0] _T_2780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5158;
  reg [31:0] _T_2781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5159;
  reg [31:0] _T_2781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5160;
  reg [31:0] _T_2782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5161;
  reg [31:0] _T_2782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5162;
  reg [31:0] _T_2783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5163;
  reg [31:0] _T_2783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5164;
  reg [31:0] _T_2784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5165;
  reg [31:0] _T_2784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5166;
  reg [31:0] _T_2785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5167;
  reg [31:0] _T_2785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5168;
  reg [31:0] _T_2786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5169;
  reg [31:0] _T_2786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5170;
  reg [31:0] _T_2787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5171;
  reg [31:0] _T_2787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5172;
  reg [31:0] _T_2788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5173;
  reg [31:0] _T_2788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5174;
  reg [31:0] _T_2789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5175;
  reg [31:0] _T_2789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5176;
  reg [31:0] _T_2790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5177;
  reg [31:0] _T_2790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5178;
  reg [31:0] _T_2791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5179;
  reg [31:0] _T_2791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5180;
  reg [31:0] _T_2792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5181;
  reg [31:0] _T_2792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5182;
  reg [31:0] _T_2793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5183;
  reg [31:0] _T_2793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5184;
  reg [31:0] _T_2794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5185;
  reg [31:0] _T_2794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5186;
  reg [31:0] _T_2795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5187;
  reg [31:0] _T_2795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5188;
  reg [31:0] _T_2796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5189;
  reg [31:0] _T_2796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5190;
  reg [31:0] _T_2797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5191;
  reg [31:0] _T_2797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5192;
  reg [31:0] _T_2798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5193;
  reg [31:0] _T_2798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5194;
  reg [31:0] _T_2799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5195;
  reg [31:0] _T_2799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5196;
  reg [31:0] _T_2800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5197;
  reg [31:0] _T_2800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5198;
  reg [31:0] _T_2801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5199;
  reg [31:0] _T_2801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5200;
  reg [31:0] _T_2802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5201;
  reg [31:0] _T_2802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5202;
  reg [31:0] _T_2803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5203;
  reg [31:0] _T_2803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5204;
  reg [31:0] _T_2804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5205;
  reg [31:0] _T_2804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5206;
  reg [31:0] _T_2805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5207;
  reg [31:0] _T_2805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5208;
  reg [31:0] _T_2806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5209;
  reg [31:0] _T_2806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5210;
  reg [31:0] _T_2807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5211;
  reg [31:0] _T_2807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5212;
  reg [31:0] _T_2808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5213;
  reg [31:0] _T_2808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5214;
  reg [31:0] _T_2809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5215;
  reg [31:0] _T_2809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5216;
  reg [31:0] _T_2810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5217;
  reg [31:0] _T_2810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5218;
  reg [31:0] _T_2811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5219;
  reg [31:0] _T_2811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5220;
  reg [31:0] _T_2812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5221;
  reg [31:0] _T_2812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5222;
  reg [31:0] _T_2813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5223;
  reg [31:0] _T_2813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5224;
  reg [31:0] _T_2814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5225;
  reg [31:0] _T_2814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5226;
  reg [31:0] _T_2815_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5227;
  reg [31:0] _T_2815_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5228;
  reg [31:0] _T_2816_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5229;
  reg [31:0] _T_2816_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5230;
  reg [31:0] _T_2817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5231;
  reg [31:0] _T_2817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5232;
  reg [31:0] _T_2818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5233;
  reg [31:0] _T_2818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5234;
  reg [31:0] _T_2819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5235;
  reg [31:0] _T_2819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5236;
  reg [31:0] _T_2820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5237;
  reg [31:0] _T_2820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5238;
  reg [31:0] _T_2821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5239;
  reg [31:0] _T_2821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5240;
  reg [31:0] _T_2822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5241;
  reg [31:0] _T_2822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5242;
  reg [31:0] _T_2823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5243;
  reg [31:0] _T_2823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5244;
  reg [31:0] _T_2824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5245;
  reg [31:0] _T_2824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5246;
  reg [31:0] _T_2825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5247;
  reg [31:0] _T_2825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5248;
  reg [31:0] _T_2826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5249;
  reg [31:0] _T_2826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5250;
  reg [31:0] _T_2827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5251;
  reg [31:0] _T_2827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5252;
  reg [31:0] _T_2828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5253;
  reg [31:0] _T_2828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5254;
  reg [31:0] _T_2829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5255;
  reg [31:0] _T_2829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5256;
  reg [31:0] _T_2830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5257;
  reg [31:0] _T_2830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5258;
  reg [31:0] _T_2831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5259;
  reg [31:0] _T_2831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5260;
  reg [31:0] _T_2832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5261;
  reg [31:0] _T_2832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5262;
  reg [31:0] _T_2833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5263;
  reg [31:0] _T_2833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5264;
  reg [31:0] _T_2834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5265;
  reg [31:0] _T_2834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5266;
  reg [31:0] _T_2835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5267;
  reg [31:0] _T_2835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5268;
  reg [31:0] _T_2836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5269;
  reg [31:0] _T_2836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5270;
  reg [31:0] _T_2837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5271;
  reg [31:0] _T_2837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5272;
  reg [31:0] _T_2838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5273;
  reg [31:0] _T_2838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5274;
  reg [31:0] _T_2839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5275;
  reg [31:0] _T_2839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5276;
  reg [31:0] _T_2840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5277;
  reg [31:0] _T_2840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5278;
  reg [31:0] _T_2841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5279;
  reg [31:0] _T_2841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5280;
  reg [31:0] _T_2842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5281;
  reg [31:0] _T_2842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5282;
  reg [31:0] _T_2843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5283;
  reg [31:0] _T_2843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5284;
  reg [31:0] _T_2844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5285;
  reg [31:0] _T_2844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5286;
  reg [31:0] _T_2845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5287;
  reg [31:0] _T_2845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5288;
  reg [31:0] _T_2846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5289;
  reg [31:0] _T_2846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5290;
  reg [31:0] _T_2847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5291;
  reg [31:0] _T_2847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5292;
  reg [31:0] _T_2848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5293;
  reg [31:0] _T_2848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5294;
  reg [31:0] _T_2849_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5295;
  reg [31:0] _T_2849_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5296;
  reg [31:0] _T_2850_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5297;
  reg [31:0] _T_2850_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5298;
  reg [31:0] _T_2851_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5299;
  reg [31:0] _T_2851_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5300;
  reg [31:0] _T_2852_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5301;
  reg [31:0] _T_2852_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5302;
  reg [31:0] _T_2853_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5303;
  reg [31:0] _T_2853_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5304;
  reg [31:0] _T_2854_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5305;
  reg [31:0] _T_2854_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5306;
  reg [31:0] _T_2855_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5307;
  reg [31:0] _T_2855_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5308;
  reg [31:0] _T_2856_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5309;
  reg [31:0] _T_2856_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5310;
  reg [31:0] _T_2857_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5311;
  reg [31:0] _T_2857_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5312;
  reg [31:0] _T_2858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5313;
  reg [31:0] _T_2858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5314;
  reg [31:0] _T_2859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5315;
  reg [31:0] _T_2859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5316;
  reg [31:0] _T_2860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5317;
  reg [31:0] _T_2860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5318;
  reg [31:0] _T_2861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5319;
  reg [31:0] _T_2861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5320;
  reg [31:0] _T_2862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5321;
  reg [31:0] _T_2862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5322;
  reg [31:0] _T_2863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5323;
  reg [31:0] _T_2863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5324;
  reg [31:0] _T_2864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5325;
  reg [31:0] _T_2864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5326;
  reg [31:0] _T_2865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5327;
  reg [31:0] _T_2865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5328;
  reg [31:0] _T_2866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5329;
  reg [31:0] _T_2866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5330;
  reg [31:0] _T_2867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5331;
  reg [31:0] _T_2867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5332;
  reg [31:0] _T_2868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5333;
  reg [31:0] _T_2868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5334;
  reg [31:0] _T_2869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5335;
  reg [31:0] _T_2869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5336;
  reg [31:0] _T_2870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5337;
  reg [31:0] _T_2870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5338;
  reg [31:0] _T_2871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5339;
  reg [31:0] _T_2871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5340;
  reg [31:0] _T_2872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5341;
  reg [31:0] _T_2872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5342;
  reg [31:0] _T_2873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5343;
  reg [31:0] _T_2873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5344;
  reg [31:0] _T_2874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5345;
  reg [31:0] _T_2874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5346;
  reg [31:0] _T_2875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5347;
  reg [31:0] _T_2875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5348;
  reg [31:0] _T_2876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5349;
  reg [31:0] _T_2876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5350;
  reg [31:0] _T_2877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5351;
  reg [31:0] _T_2877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5352;
  reg [31:0] _T_2878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5353;
  reg [31:0] _T_2878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5354;
  reg [31:0] _T_2879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5355;
  reg [31:0] _T_2879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5356;
  reg [31:0] _T_2880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5357;
  reg [31:0] _T_2880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5358;
  reg [31:0] _T_2881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5359;
  reg [31:0] _T_2881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5360;
  reg [31:0] _T_2882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5361;
  reg [31:0] _T_2882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5362;
  reg [31:0] _T_2883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5363;
  reg [31:0] _T_2883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5364;
  reg [31:0] _T_2884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5365;
  reg [31:0] _T_2884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5366;
  reg [31:0] _T_2885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5367;
  reg [31:0] _T_2885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5368;
  reg [31:0] _T_2886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5369;
  reg [31:0] _T_2886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5370;
  reg [31:0] _T_2887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5371;
  reg [31:0] _T_2887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5372;
  reg [31:0] _T_2888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5373;
  reg [31:0] _T_2888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5374;
  reg [31:0] _T_2889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5375;
  reg [31:0] _T_2889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5376;
  reg [31:0] _T_2890_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5377;
  reg [31:0] _T_2890_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5378;
  reg [31:0] _T_2891_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5379;
  reg [31:0] _T_2891_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5380;
  reg [31:0] _T_2892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5381;
  reg [31:0] _T_2892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5382;
  wire [63:0] _T_2897;
  reg [31:0] _T_2902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5383;
  reg [31:0] _T_2902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5384;
  reg [31:0] _T_2903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5385;
  reg [31:0] _T_2903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5386;
  reg [31:0] _T_2904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5387;
  reg [31:0] _T_2904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5388;
  reg [31:0] _T_2905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5389;
  reg [31:0] _T_2905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5390;
  reg [31:0] _T_2906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5391;
  reg [31:0] _T_2906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5392;
  reg [31:0] _T_2907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5393;
  reg [31:0] _T_2907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5394;
  reg [31:0] _T_2908_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5395;
  reg [31:0] _T_2908_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5396;
  reg [31:0] _T_2909_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5397;
  reg [31:0] _T_2909_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5398;
  reg [31:0] _T_2910_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5399;
  reg [31:0] _T_2910_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5400;
  reg [31:0] _T_2911_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5401;
  reg [31:0] _T_2911_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5402;
  reg [31:0] _T_2912_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5403;
  reg [31:0] _T_2912_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5404;
  reg [31:0] _T_2913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5405;
  reg [31:0] _T_2913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5406;
  reg [31:0] _T_2914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5407;
  reg [31:0] _T_2914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5408;
  reg [31:0] _T_2915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5409;
  reg [31:0] _T_2915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5410;
  reg [31:0] _T_2916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5411;
  reg [31:0] _T_2916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5412;
  reg [31:0] _T_2917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5413;
  reg [31:0] _T_2917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5414;
  reg [31:0] _T_2918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5415;
  reg [31:0] _T_2918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5416;
  reg [31:0] _T_2919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5417;
  reg [31:0] _T_2919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5418;
  reg [31:0] _T_2920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5419;
  reg [31:0] _T_2920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5420;
  reg [31:0] _T_2921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5421;
  reg [31:0] _T_2921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5422;
  reg [31:0] _T_2922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5423;
  reg [31:0] _T_2922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5424;
  reg [31:0] _T_2923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5425;
  reg [31:0] _T_2923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5426;
  reg [31:0] _T_2924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5427;
  reg [31:0] _T_2924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5428;
  reg [31:0] _T_2925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5429;
  reg [31:0] _T_2925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5430;
  reg [31:0] _T_2926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5431;
  reg [31:0] _T_2926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5432;
  reg [31:0] _T_2927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5433;
  reg [31:0] _T_2927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5434;
  reg [31:0] _T_2928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5435;
  reg [31:0] _T_2928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5436;
  reg [31:0] _T_2929_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5437;
  reg [31:0] _T_2929_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5438;
  reg [31:0] _T_2930_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5439;
  reg [31:0] _T_2930_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5440;
  reg [31:0] _T_2931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5441;
  reg [31:0] _T_2931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5442;
  reg [31:0] _T_2932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5443;
  reg [31:0] _T_2932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5444;
  reg [31:0] _T_2933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5445;
  reg [31:0] _T_2933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5446;
  reg [31:0] _T_2934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5447;
  reg [31:0] _T_2934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5448;
  reg [31:0] _T_2935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5449;
  reg [31:0] _T_2935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5450;
  reg [31:0] _T_2936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5451;
  reg [31:0] _T_2936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5452;
  reg [31:0] _T_2937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5453;
  reg [31:0] _T_2937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5454;
  reg [31:0] _T_2938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5455;
  reg [31:0] _T_2938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5456;
  reg [31:0] _T_2939_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5457;
  reg [31:0] _T_2939_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5458;
  reg [31:0] _T_2940_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5459;
  reg [31:0] _T_2940_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5460;
  reg [31:0] _T_2941_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5461;
  reg [31:0] _T_2941_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5462;
  reg [31:0] _T_2942_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5463;
  reg [31:0] _T_2942_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5464;
  reg [31:0] _T_2943_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5465;
  reg [31:0] _T_2943_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5466;
  reg [31:0] _T_2944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5467;
  reg [31:0] _T_2944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5468;
  reg [31:0] _T_2945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5469;
  reg [31:0] _T_2945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5470;
  reg [31:0] _T_2946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5471;
  reg [31:0] _T_2946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5472;
  reg [31:0] _T_2947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5473;
  reg [31:0] _T_2947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5474;
  reg [31:0] _T_2948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5475;
  reg [31:0] _T_2948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5476;
  reg [31:0] _T_2949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5477;
  reg [31:0] _T_2949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5478;
  reg [31:0] _T_2950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5479;
  reg [31:0] _T_2950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5480;
  reg [31:0] _T_2951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5481;
  reg [31:0] _T_2951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5482;
  reg [31:0] _T_2952_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5483;
  reg [31:0] _T_2952_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5484;
  reg [31:0] _T_2953_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5485;
  reg [31:0] _T_2953_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5486;
  reg [31:0] _T_2954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5487;
  reg [31:0] _T_2954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5488;
  reg [31:0] _T_2955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5489;
  reg [31:0] _T_2955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5490;
  reg [31:0] _T_2956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5491;
  reg [31:0] _T_2956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5492;
  reg [31:0] _T_2957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5493;
  reg [31:0] _T_2957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5494;
  reg [31:0] _T_2958_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5495;
  reg [31:0] _T_2958_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5496;
  reg [31:0] _T_2959_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5497;
  reg [31:0] _T_2959_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5498;
  reg [31:0] _T_2960_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5499;
  reg [31:0] _T_2960_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5500;
  reg [31:0] _T_2961_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5501;
  reg [31:0] _T_2961_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5502;
  reg [31:0] _T_2962_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5503;
  reg [31:0] _T_2962_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5504;
  reg [31:0] _T_2963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5505;
  reg [31:0] _T_2963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5506;
  reg [31:0] _T_2964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5507;
  reg [31:0] _T_2964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5508;
  reg [31:0] _T_2965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5509;
  reg [31:0] _T_2965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5510;
  reg [31:0] _T_2966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5511;
  reg [31:0] _T_2966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5512;
  reg [31:0] _T_2967_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5513;
  reg [31:0] _T_2967_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5514;
  reg [31:0] _T_2968_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5515;
  reg [31:0] _T_2968_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5516;
  reg [31:0] _T_2969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5517;
  reg [31:0] _T_2969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5518;
  reg [31:0] _T_2970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5519;
  reg [31:0] _T_2970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5520;
  reg [31:0] _T_2971_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5521;
  reg [31:0] _T_2971_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5522;
  reg [31:0] _T_2972_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5523;
  reg [31:0] _T_2972_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5524;
  reg [31:0] _T_2973_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5525;
  reg [31:0] _T_2973_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5526;
  reg [31:0] _T_2974_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5527;
  reg [31:0] _T_2974_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5528;
  reg [31:0] _T_2975_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5529;
  reg [31:0] _T_2975_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5530;
  reg [31:0] _T_2976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5531;
  reg [31:0] _T_2976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5532;
  reg [31:0] _T_2977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5533;
  reg [31:0] _T_2977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5534;
  reg [31:0] _T_2978_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5535;
  reg [31:0] _T_2978_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5536;
  reg [31:0] _T_2979_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5537;
  reg [31:0] _T_2979_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5538;
  reg [31:0] _T_2980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5539;
  reg [31:0] _T_2980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5540;
  reg [31:0] _T_2981_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5541;
  reg [31:0] _T_2981_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5542;
  reg [31:0] _T_2982_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5543;
  reg [31:0] _T_2982_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5544;
  reg [31:0] _T_2983_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5545;
  reg [31:0] _T_2983_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5546;
  reg [31:0] _T_2984_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5547;
  reg [31:0] _T_2984_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5548;
  reg [31:0] _T_2985_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5549;
  reg [31:0] _T_2985_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5550;
  reg [31:0] _T_2986_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5551;
  reg [31:0] _T_2986_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5552;
  reg [31:0] _T_2987_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5553;
  reg [31:0] _T_2987_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5554;
  reg [31:0] _T_2988_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5555;
  reg [31:0] _T_2988_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5556;
  reg [31:0] _T_2989_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5557;
  reg [31:0] _T_2989_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5558;
  reg [31:0] _T_2990_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5559;
  reg [31:0] _T_2990_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5560;
  reg [31:0] _T_2991_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5561;
  reg [31:0] _T_2991_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5562;
  reg [31:0] _T_2992_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5563;
  reg [31:0] _T_2992_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5564;
  reg [31:0] _T_2993_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5565;
  reg [31:0] _T_2993_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5566;
  reg [31:0] _T_2994_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5567;
  reg [31:0] _T_2994_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5568;
  reg [31:0] _T_2995_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5569;
  reg [31:0] _T_2995_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5570;
  reg [31:0] _T_2996_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5571;
  reg [31:0] _T_2996_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5572;
  reg [31:0] _T_2997_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5573;
  reg [31:0] _T_2997_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5574;
  reg [31:0] _T_2998_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5575;
  reg [31:0] _T_2998_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5576;
  reg [31:0] _T_2999_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5577;
  reg [31:0] _T_2999_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5578;
  reg [31:0] _T_3000_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5579;
  reg [31:0] _T_3000_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5580;
  reg [31:0] _T_3001_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5581;
  reg [31:0] _T_3001_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5582;
  reg [31:0] _T_3002_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5583;
  reg [31:0] _T_3002_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5584;
  reg [31:0] _T_3003_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5585;
  reg [31:0] _T_3003_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5586;
  reg [31:0] _T_3004_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5587;
  reg [31:0] _T_3004_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5588;
  reg [31:0] _T_3005_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5589;
  reg [31:0] _T_3005_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5590;
  reg [31:0] _T_3006_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5591;
  reg [31:0] _T_3006_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5592;
  reg [31:0] _T_3007_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5593;
  reg [31:0] _T_3007_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5594;
  reg [31:0] _T_3008_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5595;
  reg [31:0] _T_3008_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5596;
  reg [31:0] _T_3009_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5597;
  reg [31:0] _T_3009_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5598;
  reg [31:0] _T_3010_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5599;
  reg [31:0] _T_3010_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5600;
  reg [31:0] _T_3011_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5601;
  reg [31:0] _T_3011_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5602;
  reg [31:0] _T_3012_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5603;
  reg [31:0] _T_3012_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5604;
  reg [31:0] _T_3013_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5605;
  reg [31:0] _T_3013_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5606;
  reg [31:0] _T_3014_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5607;
  reg [31:0] _T_3014_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5608;
  reg [31:0] _T_3015_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5609;
  reg [31:0] _T_3015_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5610;
  reg [31:0] _T_3016_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5611;
  reg [31:0] _T_3016_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5612;
  reg [31:0] _T_3017_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5613;
  reg [31:0] _T_3017_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5614;
  reg [31:0] _T_3018_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5615;
  reg [31:0] _T_3018_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5616;
  reg [31:0] _T_3019_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5617;
  reg [31:0] _T_3019_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5618;
  reg [31:0] _T_3020_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5619;
  reg [31:0] _T_3020_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5620;
  reg [31:0] _T_3021_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5621;
  reg [31:0] _T_3021_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5622;
  reg [31:0] _T_3022_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5623;
  reg [31:0] _T_3022_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5624;
  reg [31:0] _T_3023_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5625;
  reg [31:0] _T_3023_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5626;
  reg [31:0] _T_3024_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5627;
  reg [31:0] _T_3024_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5628;
  reg [31:0] _T_3025_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5629;
  reg [31:0] _T_3025_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5630;
  reg [31:0] _T_3026_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5631;
  reg [31:0] _T_3026_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5632;
  reg [31:0] _T_3027_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5633;
  reg [31:0] _T_3027_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5634;
  reg [31:0] _T_3028_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5635;
  reg [31:0] _T_3028_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5636;
  reg [31:0] _T_3029_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5637;
  reg [31:0] _T_3029_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5638;
  reg [31:0] _T_3032_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5639;
  reg [31:0] _T_3032_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5640;
  reg [31:0] _T_3033_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5641;
  reg [31:0] _T_3033_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5642;
  reg [31:0] _T_3034_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5643;
  reg [31:0] _T_3034_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5644;
  reg [31:0] _T_3035_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5645;
  reg [31:0] _T_3035_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5646;
  reg [31:0] _T_3036_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5647;
  reg [31:0] _T_3036_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5648;
  reg [31:0] _T_3037_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5649;
  reg [31:0] _T_3037_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5650;
  reg [31:0] _T_3038_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5651;
  reg [31:0] _T_3038_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5652;
  reg [31:0] _T_3039_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5653;
  reg [31:0] _T_3039_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5654;
  reg [31:0] _T_3040_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5655;
  reg [31:0] _T_3040_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5656;
  reg [31:0] _T_3041_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5657;
  reg [31:0] _T_3041_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5658;
  reg [31:0] _T_3042_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5659;
  reg [31:0] _T_3042_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5660;
  reg [31:0] _T_3043_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5661;
  reg [31:0] _T_3043_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5662;
  reg [31:0] _T_3044_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5663;
  reg [31:0] _T_3044_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5664;
  reg [31:0] _T_3045_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5665;
  reg [31:0] _T_3045_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5666;
  reg [31:0] _T_3046_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5667;
  reg [31:0] _T_3046_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5668;
  reg [31:0] _T_3047_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5669;
  reg [31:0] _T_3047_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5670;
  reg [31:0] _T_3048_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5671;
  reg [31:0] _T_3048_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5672;
  reg [31:0] _T_3049_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5673;
  reg [31:0] _T_3049_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5674;
  reg [31:0] _T_3050_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5675;
  reg [31:0] _T_3050_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5676;
  reg [31:0] _T_3051_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5677;
  reg [31:0] _T_3051_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5678;
  reg [31:0] _T_3052_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5679;
  reg [31:0] _T_3052_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5680;
  reg [31:0] _T_3053_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5681;
  reg [31:0] _T_3053_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5682;
  reg [31:0] _T_3054_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5683;
  reg [31:0] _T_3054_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5684;
  reg [31:0] _T_3055_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5685;
  reg [31:0] _T_3055_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5686;
  reg [31:0] _T_3056_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5687;
  reg [31:0] _T_3056_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5688;
  reg [31:0] _T_3057_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5689;
  reg [31:0] _T_3057_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5690;
  reg [31:0] _T_3058_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5691;
  reg [31:0] _T_3058_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5692;
  reg [31:0] _T_3059_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5693;
  reg [31:0] _T_3059_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5694;
  reg [31:0] _T_3060_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5695;
  reg [31:0] _T_3060_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5696;
  reg [31:0] _T_3061_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5697;
  reg [31:0] _T_3061_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5698;
  reg [31:0] _T_3062_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5699;
  reg [31:0] _T_3062_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5700;
  reg [31:0] _T_3063_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5701;
  reg [31:0] _T_3063_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5702;
  reg [31:0] _T_3064_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5703;
  reg [31:0] _T_3064_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5704;
  reg [31:0] _T_3065_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5705;
  reg [31:0] _T_3065_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5706;
  reg [31:0] _T_3066_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5707;
  reg [31:0] _T_3066_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5708;
  reg [31:0] _T_3067_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5709;
  reg [31:0] _T_3067_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5710;
  reg [31:0] _T_3068_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5711;
  reg [31:0] _T_3068_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5712;
  reg [31:0] _T_3069_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5713;
  reg [31:0] _T_3069_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5714;
  reg [31:0] _T_3070_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5715;
  reg [31:0] _T_3070_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5716;
  reg [31:0] _T_3071_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5717;
  reg [31:0] _T_3071_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5718;
  reg [31:0] _T_3072_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5719;
  reg [31:0] _T_3072_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5720;
  reg [31:0] _T_3073_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5721;
  reg [31:0] _T_3073_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5722;
  reg [31:0] _T_3074_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5723;
  reg [31:0] _T_3074_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5724;
  reg [31:0] _T_3075_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5725;
  reg [31:0] _T_3075_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5726;
  reg [31:0] _T_3076_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5727;
  reg [31:0] _T_3076_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5728;
  reg [31:0] _T_3077_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5729;
  reg [31:0] _T_3077_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5730;
  reg [31:0] _T_3078_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5731;
  reg [31:0] _T_3078_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5732;
  reg [31:0] _T_3079_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5733;
  reg [31:0] _T_3079_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5734;
  reg [31:0] _T_3080_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5735;
  reg [31:0] _T_3080_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5736;
  reg [31:0] _T_3081_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5737;
  reg [31:0] _T_3081_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5738;
  reg [31:0] _T_3082_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5739;
  reg [31:0] _T_3082_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5740;
  reg [31:0] _T_3083_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5741;
  reg [31:0] _T_3083_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5742;
  reg [31:0] _T_3084_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5743;
  reg [31:0] _T_3084_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5744;
  reg [31:0] _T_3085_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5745;
  reg [31:0] _T_3085_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5746;
  reg [31:0] _T_3086_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5747;
  reg [31:0] _T_3086_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5748;
  reg [31:0] _T_3087_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5749;
  reg [31:0] _T_3087_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5750;
  reg [31:0] _T_3088_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5751;
  reg [31:0] _T_3088_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5752;
  reg [31:0] _T_3089_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5753;
  reg [31:0] _T_3089_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5754;
  reg [31:0] _T_3090_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5755;
  reg [31:0] _T_3090_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5756;
  reg [31:0] _T_3091_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5757;
  reg [31:0] _T_3091_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5758;
  reg [31:0] _T_3092_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5759;
  reg [31:0] _T_3092_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5760;
  reg [31:0] _T_3093_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5761;
  reg [31:0] _T_3093_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5762;
  reg [31:0] _T_3094_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5763;
  reg [31:0] _T_3094_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5764;
  reg [31:0] _T_3095_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5765;
  reg [31:0] _T_3095_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5766;
  wire [63:0] _T_3100;
  reg [31:0] _T_3105_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5767;
  reg [31:0] _T_3105_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5768;
  reg [31:0] _T_3106_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5769;
  reg [31:0] _T_3106_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5770;
  reg [31:0] _T_3107_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5771;
  reg [31:0] _T_3107_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5772;
  reg [31:0] _T_3108_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5773;
  reg [31:0] _T_3108_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5774;
  reg [31:0] _T_3109_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5775;
  reg [31:0] _T_3109_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5776;
  reg [31:0] _T_3110_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5777;
  reg [31:0] _T_3110_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5778;
  reg [31:0] _T_3111_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5779;
  reg [31:0] _T_3111_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5780;
  reg [31:0] _T_3112_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5781;
  reg [31:0] _T_3112_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5782;
  reg [31:0] _T_3113_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5783;
  reg [31:0] _T_3113_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5784;
  reg [31:0] _T_3114_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5785;
  reg [31:0] _T_3114_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5786;
  reg [31:0] _T_3115_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5787;
  reg [31:0] _T_3115_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5788;
  reg [31:0] _T_3116_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5789;
  reg [31:0] _T_3116_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5790;
  reg [31:0] _T_3117_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5791;
  reg [31:0] _T_3117_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5792;
  reg [31:0] _T_3118_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5793;
  reg [31:0] _T_3118_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5794;
  reg [31:0] _T_3119_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5795;
  reg [31:0] _T_3119_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5796;
  reg [31:0] _T_3120_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5797;
  reg [31:0] _T_3120_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5798;
  reg [31:0] _T_3121_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5799;
  reg [31:0] _T_3121_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5800;
  reg [31:0] _T_3122_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5801;
  reg [31:0] _T_3122_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5802;
  reg [31:0] _T_3123_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5803;
  reg [31:0] _T_3123_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5804;
  reg [31:0] _T_3124_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5805;
  reg [31:0] _T_3124_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5806;
  reg [31:0] _T_3125_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5807;
  reg [31:0] _T_3125_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5808;
  reg [31:0] _T_3126_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5809;
  reg [31:0] _T_3126_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5810;
  reg [31:0] _T_3127_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5811;
  reg [31:0] _T_3127_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5812;
  reg [31:0] _T_3128_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5813;
  reg [31:0] _T_3128_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5814;
  reg [31:0] _T_3129_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5815;
  reg [31:0] _T_3129_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5816;
  reg [31:0] _T_3130_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5817;
  reg [31:0] _T_3130_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5818;
  reg [31:0] _T_3131_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5819;
  reg [31:0] _T_3131_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5820;
  reg [31:0] _T_3132_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5821;
  reg [31:0] _T_3132_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5822;
  reg [31:0] _T_3133_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5823;
  reg [31:0] _T_3133_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5824;
  reg [31:0] _T_3134_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5825;
  reg [31:0] _T_3134_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5826;
  reg [31:0] _T_3135_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5827;
  reg [31:0] _T_3135_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5828;
  reg [31:0] _T_3136_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5829;
  reg [31:0] _T_3136_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5830;
  reg [31:0] _T_3137_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5831;
  reg [31:0] _T_3137_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5832;
  reg [31:0] _T_3138_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5833;
  reg [31:0] _T_3138_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5834;
  reg [31:0] _T_3139_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5835;
  reg [31:0] _T_3139_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5836;
  reg [31:0] _T_3140_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5837;
  reg [31:0] _T_3140_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5838;
  reg [31:0] _T_3141_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5839;
  reg [31:0] _T_3141_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5840;
  reg [31:0] _T_3142_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5841;
  reg [31:0] _T_3142_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5842;
  reg [31:0] _T_3143_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5843;
  reg [31:0] _T_3143_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5844;
  reg [31:0] _T_3144_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5845;
  reg [31:0] _T_3144_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5846;
  reg [31:0] _T_3145_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5847;
  reg [31:0] _T_3145_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5848;
  reg [31:0] _T_3146_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5849;
  reg [31:0] _T_3146_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5850;
  reg [31:0] _T_3147_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5851;
  reg [31:0] _T_3147_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5852;
  reg [31:0] _T_3148_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5853;
  reg [31:0] _T_3148_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5854;
  reg [31:0] _T_3149_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5855;
  reg [31:0] _T_3149_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5856;
  reg [31:0] _T_3150_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5857;
  reg [31:0] _T_3150_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5858;
  reg [31:0] _T_3151_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5859;
  reg [31:0] _T_3151_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5860;
  reg [31:0] _T_3152_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5861;
  reg [31:0] _T_3152_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5862;
  reg [31:0] _T_3153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5863;
  reg [31:0] _T_3153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5864;
  reg [31:0] _T_3154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5865;
  reg [31:0] _T_3154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5866;
  reg [31:0] _T_3155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5867;
  reg [31:0] _T_3155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5868;
  reg [31:0] _T_3156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5869;
  reg [31:0] _T_3156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5870;
  reg [31:0] _T_3157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5871;
  reg [31:0] _T_3157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5872;
  reg [31:0] _T_3158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5873;
  reg [31:0] _T_3158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5874;
  reg [31:0] _T_3159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5875;
  reg [31:0] _T_3159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5876;
  reg [31:0] _T_3160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5877;
  reg [31:0] _T_3160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5878;
  reg [31:0] _T_3161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5879;
  reg [31:0] _T_3161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5880;
  reg [31:0] _T_3162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5881;
  reg [31:0] _T_3162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5882;
  reg [31:0] _T_3163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5883;
  reg [31:0] _T_3163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5884;
  reg [31:0] _T_3164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5885;
  reg [31:0] _T_3164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5886;
  reg [31:0] _T_3165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5887;
  reg [31:0] _T_3165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5888;
  reg [31:0] _T_3166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5889;
  reg [31:0] _T_3166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5890;
  reg [31:0] _T_3167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5891;
  reg [31:0] _T_3167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5892;
  reg [31:0] _T_3168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5893;
  reg [31:0] _T_3168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5894;
  reg [31:0] _T_3171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5895;
  reg [31:0] _T_3171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5896;
  reg [31:0] _T_3172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5897;
  reg [31:0] _T_3172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5898;
  reg [31:0] _T_3173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5899;
  reg [31:0] _T_3173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5900;
  reg [31:0] _T_3174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5901;
  reg [31:0] _T_3174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5902;
  reg [31:0] _T_3175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5903;
  reg [31:0] _T_3175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5904;
  reg [31:0] _T_3176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5905;
  reg [31:0] _T_3176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5906;
  reg [31:0] _T_3177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5907;
  reg [31:0] _T_3177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5908;
  reg [31:0] _T_3178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5909;
  reg [31:0] _T_3178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5910;
  reg [31:0] _T_3179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5911;
  reg [31:0] _T_3179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5912;
  reg [31:0] _T_3180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5913;
  reg [31:0] _T_3180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5914;
  reg [31:0] _T_3181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5915;
  reg [31:0] _T_3181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5916;
  reg [31:0] _T_3182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5917;
  reg [31:0] _T_3182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5918;
  reg [31:0] _T_3183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5919;
  reg [31:0] _T_3183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5920;
  reg [31:0] _T_3184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5921;
  reg [31:0] _T_3184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5922;
  reg [31:0] _T_3185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5923;
  reg [31:0] _T_3185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5924;
  reg [31:0] _T_3186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5925;
  reg [31:0] _T_3186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5926;
  reg [31:0] _T_3187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5927;
  reg [31:0] _T_3187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5928;
  reg [31:0] _T_3188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5929;
  reg [31:0] _T_3188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5930;
  reg [31:0] _T_3189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5931;
  reg [31:0] _T_3189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5932;
  reg [31:0] _T_3190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5933;
  reg [31:0] _T_3190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5934;
  reg [31:0] _T_3191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5935;
  reg [31:0] _T_3191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5936;
  reg [31:0] _T_3192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5937;
  reg [31:0] _T_3192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5938;
  reg [31:0] _T_3193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5939;
  reg [31:0] _T_3193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5940;
  reg [31:0] _T_3194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5941;
  reg [31:0] _T_3194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5942;
  reg [31:0] _T_3195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5943;
  reg [31:0] _T_3195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5944;
  reg [31:0] _T_3196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5945;
  reg [31:0] _T_3196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5946;
  reg [31:0] _T_3197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5947;
  reg [31:0] _T_3197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5948;
  reg [31:0] _T_3198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5949;
  reg [31:0] _T_3198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5950;
  reg [31:0] _T_3199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5951;
  reg [31:0] _T_3199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5952;
  reg [31:0] _T_3200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5953;
  reg [31:0] _T_3200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5954;
  reg [31:0] _T_3201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5955;
  reg [31:0] _T_3201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5956;
  reg [31:0] _T_3202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5957;
  reg [31:0] _T_3202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5958;
  wire [63:0] _T_3207;
  reg [31:0] _T_3212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5959;
  reg [31:0] _T_3212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5960;
  reg [31:0] _T_3213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5961;
  reg [31:0] _T_3213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5962;
  reg [31:0] _T_3214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5963;
  reg [31:0] _T_3214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5964;
  reg [31:0] _T_3215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5965;
  reg [31:0] _T_3215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5966;
  reg [31:0] _T_3216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5967;
  reg [31:0] _T_3216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5968;
  reg [31:0] _T_3217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5969;
  reg [31:0] _T_3217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5970;
  reg [31:0] _T_3218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5971;
  reg [31:0] _T_3218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5972;
  reg [31:0] _T_3219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5973;
  reg [31:0] _T_3219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5974;
  reg [31:0] _T_3220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5975;
  reg [31:0] _T_3220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5976;
  reg [31:0] _T_3221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5977;
  reg [31:0] _T_3221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5978;
  reg [31:0] _T_3222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5979;
  reg [31:0] _T_3222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5980;
  reg [31:0] _T_3223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5981;
  reg [31:0] _T_3223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5982;
  reg [31:0] _T_3224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5983;
  reg [31:0] _T_3224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5984;
  reg [31:0] _T_3225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5985;
  reg [31:0] _T_3225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5986;
  reg [31:0] _T_3226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5987;
  reg [31:0] _T_3226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5988;
  reg [31:0] _T_3227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5989;
  reg [31:0] _T_3227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5990;
  reg [31:0] _T_3228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5991;
  reg [31:0] _T_3228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5992;
  reg [31:0] _T_3229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5993;
  reg [31:0] _T_3229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5994;
  reg [31:0] _T_3230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5995;
  reg [31:0] _T_3230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5996;
  reg [31:0] _T_3231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5997;
  reg [31:0] _T_3231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5998;
  reg [31:0] _T_3232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5999;
  reg [31:0] _T_3232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6000;
  reg [31:0] _T_3233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6001;
  reg [31:0] _T_3233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6002;
  reg [31:0] _T_3234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6003;
  reg [31:0] _T_3234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6004;
  reg [31:0] _T_3235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6005;
  reg [31:0] _T_3235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6006;
  reg [31:0] _T_3236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6007;
  reg [31:0] _T_3236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6008;
  reg [31:0] _T_3237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6009;
  reg [31:0] _T_3237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6010;
  reg [31:0] _T_3238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6011;
  reg [31:0] _T_3238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6012;
  reg [31:0] _T_3239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6013;
  reg [31:0] _T_3239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6014;
  reg [31:0] _T_3240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6015;
  reg [31:0] _T_3240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6016;
  reg [31:0] _T_3241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6017;
  reg [31:0] _T_3241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6018;
  reg [31:0] _T_3242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6019;
  reg [31:0] _T_3242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6020;
  reg [31:0] _T_3243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6021;
  reg [31:0] _T_3243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6022;
  reg [31:0] _T_3246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6023;
  reg [31:0] _T_3246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6024;
  reg [31:0] _T_3247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6025;
  reg [31:0] _T_3247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6026;
  reg [31:0] _T_3248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6027;
  reg [31:0] _T_3248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6028;
  reg [31:0] _T_3249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6029;
  reg [31:0] _T_3249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6030;
  reg [31:0] _T_3250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6031;
  reg [31:0] _T_3250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6032;
  reg [31:0] _T_3251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6033;
  reg [31:0] _T_3251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6034;
  reg [31:0] _T_3252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6035;
  reg [31:0] _T_3252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6036;
  reg [31:0] _T_3253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6037;
  reg [31:0] _T_3253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6038;
  reg [31:0] _T_3254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6039;
  reg [31:0] _T_3254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6040;
  reg [31:0] _T_3255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6041;
  reg [31:0] _T_3255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6042;
  reg [31:0] _T_3256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6043;
  reg [31:0] _T_3256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6044;
  reg [31:0] _T_3257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6045;
  reg [31:0] _T_3257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6046;
  reg [31:0] _T_3258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6047;
  reg [31:0] _T_3258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6048;
  reg [31:0] _T_3259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6049;
  reg [31:0] _T_3259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6050;
  reg [31:0] _T_3260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6051;
  reg [31:0] _T_3260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6052;
  reg [31:0] _T_3261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6053;
  reg [31:0] _T_3261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6054;
  wire [31:0] _GEN_6050; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6051; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6052; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6053; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6054; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6055; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6056; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6057; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6058; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6059; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6060; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6061; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6062; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6063; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6066; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6067; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6068; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6069; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6070; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6071; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6072; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6073; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6074; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6075; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6076; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6077; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6078; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6079; // @[FFT.scala 35:12]
  reg [31:0] _T_3267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6055;
  reg [31:0] _T_3267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6056;
  reg [31:0] _T_3268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6057;
  reg [31:0] _T_3268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6058;
  reg [31:0] _T_3269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6059;
  reg [31:0] _T_3269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6060;
  reg [31:0] _T_3270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6061;
  reg [31:0] _T_3270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6062;
  reg [31:0] _T_3271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6063;
  reg [31:0] _T_3271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6064;
  reg [31:0] _T_3272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6065;
  reg [31:0] _T_3272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6066;
  reg [31:0] _T_3273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6067;
  reg [31:0] _T_3273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6068;
  reg [31:0] _T_3274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6069;
  reg [31:0] _T_3274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6070;
  reg [31:0] _T_3275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6071;
  reg [31:0] _T_3275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6072;
  reg [31:0] _T_3276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6073;
  reg [31:0] _T_3276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6074;
  reg [31:0] _T_3277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6075;
  reg [31:0] _T_3277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6076;
  reg [31:0] _T_3278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6077;
  reg [31:0] _T_3278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6078;
  reg [31:0] _T_3279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6079;
  reg [31:0] _T_3279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6080;
  reg [31:0] _T_3280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6081;
  reg [31:0] _T_3280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6082;
  reg [31:0] _T_3281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6083;
  reg [31:0] _T_3281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6084;
  reg [31:0] _T_3282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6085;
  reg [31:0] _T_3282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6086;
  reg [31:0] _T_3285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6087;
  reg [31:0] _T_3285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6088;
  reg [31:0] _T_3286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6089;
  reg [31:0] _T_3286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6090;
  reg [31:0] _T_3287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6091;
  reg [31:0] _T_3287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6092;
  reg [31:0] _T_3288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6093;
  reg [31:0] _T_3288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6094;
  reg [31:0] _T_3289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6095;
  reg [31:0] _T_3289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6096;
  reg [31:0] _T_3290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6097;
  reg [31:0] _T_3290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6098;
  reg [31:0] _T_3291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6099;
  reg [31:0] _T_3291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6100;
  reg [31:0] _T_3292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6101;
  reg [31:0] _T_3292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6102;
  wire [31:0] _GEN_6130; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6131; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6132; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6133; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6134; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6135; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6138; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6139; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6140; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6141; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6142; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6143; // @[FFT.scala 35:12]
  reg [31:0] _T_3298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6103;
  reg [31:0] _T_3298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6104;
  reg [31:0] _T_3299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6105;
  reg [31:0] _T_3299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6106;
  reg [31:0] _T_3300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6107;
  reg [31:0] _T_3300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6108;
  reg [31:0] _T_3301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6109;
  reg [31:0] _T_3301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6110;
  reg [31:0] _T_3302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6111;
  reg [31:0] _T_3302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6112;
  reg [31:0] _T_3303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6113;
  reg [31:0] _T_3303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6114;
  reg [31:0] _T_3304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6115;
  reg [31:0] _T_3304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6116;
  reg [31:0] _T_3305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6117;
  reg [31:0] _T_3305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6118;
  reg [31:0] _T_3308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6119;
  reg [31:0] _T_3308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6120;
  reg [31:0] _T_3309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6121;
  reg [31:0] _T_3309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6122;
  reg [31:0] _T_3310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6123;
  reg [31:0] _T_3310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6124;
  reg [31:0] _T_3311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6125;
  reg [31:0] _T_3311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6126;
  wire [31:0] _GEN_6170; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6171; // @[FFT.scala 34:12]
  wire [31:0] _GEN_6174; // @[FFT.scala 35:12]
  wire [31:0] _GEN_6175; // @[FFT.scala 35:12]
  reg [31:0] _T_3317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6127;
  reg [31:0] _T_3317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6128;
  reg [31:0] _T_3318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6129;
  reg [31:0] _T_3318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6130;
  reg [31:0] _T_3319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6131;
  reg [31:0] _T_3319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6132;
  reg [31:0] _T_3320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6133;
  reg [31:0] _T_3320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6134;
  reg [31:0] _T_3323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6135;
  reg [31:0] _T_3323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6136;
  reg [31:0] _T_3324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6137;
  reg [31:0] _T_3324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6138;
  reg [31:0] _T_3330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6139;
  reg [31:0] _T_3330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6140;
  reg [31:0] _T_3331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6141;
  reg [31:0] _T_3331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6142;
  reg [31:0] _T_3334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6143;
  reg [31:0] _T_3334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6144;
  reg [31:0] out1D1_re; // @[FFT.scala 81:23]
  reg [31:0] _RAND_6145;
  reg [31:0] out1D1_im; // @[FFT.scala 81:23]
  reg [31:0] _RAND_6146;
  reg [31:0] _T_3335_re; // @[FFT.scala 85:22]
  reg [31:0] _RAND_6147;
  reg [31:0] _T_3335_im; // @[FFT.scala 85:22]
  reg [31:0] _RAND_6148;
  reg [31:0] _T_3336_re; // @[FFT.scala 86:22]
  reg [31:0] _RAND_6149;
  reg [31:0] _T_3336_im; // @[FFT.scala 86:22]
  reg [31:0] _RAND_6150;
  BRAM #(.ADDR_WIDTH(10), .DATA_WIDTH(64)) BRAM ( // @[FFT.scala 62:23]
    .clock(BRAM_clock),
    .en(BRAM_en),
    .addr(BRAM_addr),
    .dout(BRAM_dout)
  );
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(9), .DATA_WIDTH(64)) BRAM_1 ( // @[FFT.scala 62:23]
    .clock(BRAM_1_clock),
    .en(BRAM_1_en),
    .addr(BRAM_1_addr),
    .dout(BRAM_1_dout)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(8), .DATA_WIDTH(64)) BRAM_2 ( // @[FFT.scala 62:23]
    .clock(BRAM_2_clock),
    .en(BRAM_2_en),
    .addr(BRAM_2_addr),
    .dout(BRAM_2_dout)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(7), .DATA_WIDTH(64)) BRAM_3 ( // @[FFT.scala 62:23]
    .clock(BRAM_3_clock),
    .en(BRAM_3_en),
    .addr(BRAM_3_addr),
    .dout(BRAM_3_dout)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(6), .DATA_WIDTH(64)) BRAM_4 ( // @[FFT.scala 62:23]
    .clock(BRAM_4_clock),
    .en(BRAM_4_en),
    .addr(BRAM_4_addr),
    .dout(BRAM_4_dout)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(5), .DATA_WIDTH(64)) BRAM_5 ( // @[FFT.scala 62:23]
    .clock(BRAM_5_clock),
    .en(BRAM_5_en),
    .addr(BRAM_5_addr),
    .dout(BRAM_5_dout)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  Butterfly Butterfly_8 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_8_io_in1_re),
    .io_in1_im(Butterfly_8_io_in1_im),
    .io_in2_re(Butterfly_8_io_in2_re),
    .io_in2_im(Butterfly_8_io_in2_im),
    .io_wn_re(Butterfly_8_io_wn_re),
    .io_wn_im(Butterfly_8_io_wn_im),
    .io_out1_re(Butterfly_8_io_out1_re),
    .io_out1_im(Butterfly_8_io_out1_im),
    .io_out2_re(Butterfly_8_io_out2_re),
    .io_out2_im(Butterfly_8_io_out2_im)
  );
  Switch Switch_8 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_8_io_in1_re),
    .io_in1_im(Switch_8_io_in1_im),
    .io_in2_re(Switch_8_io_in2_re),
    .io_in2_im(Switch_8_io_in2_im),
    .io_sel(Switch_8_io_sel),
    .io_out1_re(Switch_8_io_out1_re),
    .io_out1_im(Switch_8_io_out1_im),
    .io_out2_re(Switch_8_io_out2_re),
    .io_out2_im(Switch_8_io_out2_im)
  );
  Butterfly Butterfly_9 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_9_io_in1_re),
    .io_in1_im(Butterfly_9_io_in1_im),
    .io_in2_re(Butterfly_9_io_in2_re),
    .io_in2_im(Butterfly_9_io_in2_im),
    .io_wn_re(Butterfly_9_io_wn_re),
    .io_wn_im(Butterfly_9_io_wn_im),
    .io_out1_re(Butterfly_9_io_out1_re),
    .io_out1_im(Butterfly_9_io_out1_im),
    .io_out2_re(Butterfly_9_io_out2_re),
    .io_out2_im(Butterfly_9_io_out2_im)
  );
  Switch Switch_9 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_9_io_in1_re),
    .io_in1_im(Switch_9_io_in1_im),
    .io_in2_re(Switch_9_io_in2_re),
    .io_in2_im(Switch_9_io_in2_im),
    .io_sel(Switch_9_io_sel),
    .io_out1_re(Switch_9_io_out1_re),
    .io_out1_im(Switch_9_io_out1_im),
    .io_out2_re(Switch_9_io_out2_re),
    .io_out2_im(Switch_9_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign _T_1 = cnt + 11'h1; // @[FFT.scala 42:16]
  assign _T_176 = BRAM_dout;
  assign _T_1723 = BRAM_1_dout;
  assign _T_2502 = BRAM_2_dout;
  assign _T_2897 = BRAM_3_dout;
  assign _T_3100 = BRAM_4_dout;
  assign _T_3207 = BRAM_5_dout;
  assign _GEN_6050 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_6051 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_6050); // @[FFT.scala 34:12]
  assign _GEN_6052 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_6051); // @[FFT.scala 34:12]
  assign _GEN_6053 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_6052); // @[FFT.scala 34:12]
  assign _GEN_6054 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_6053); // @[FFT.scala 34:12]
  assign _GEN_6055 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_6054); // @[FFT.scala 34:12]
  assign _GEN_6056 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_6055); // @[FFT.scala 34:12]
  assign _GEN_6057 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_6056); // @[FFT.scala 34:12]
  assign _GEN_6058 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_6057); // @[FFT.scala 34:12]
  assign _GEN_6059 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_6058); // @[FFT.scala 34:12]
  assign _GEN_6060 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_6059); // @[FFT.scala 34:12]
  assign _GEN_6061 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_6060); // @[FFT.scala 34:12]
  assign _GEN_6062 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_6061); // @[FFT.scala 34:12]
  assign _GEN_6063 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_6062); // @[FFT.scala 34:12]
  assign _GEN_6066 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_6067 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_6066); // @[FFT.scala 35:12]
  assign _GEN_6068 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_6067); // @[FFT.scala 35:12]
  assign _GEN_6069 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_6068); // @[FFT.scala 35:12]
  assign _GEN_6070 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_6069); // @[FFT.scala 35:12]
  assign _GEN_6071 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_6070); // @[FFT.scala 35:12]
  assign _GEN_6072 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_6071); // @[FFT.scala 35:12]
  assign _GEN_6073 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_6072); // @[FFT.scala 35:12]
  assign _GEN_6074 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_6073); // @[FFT.scala 35:12]
  assign _GEN_6075 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_6074); // @[FFT.scala 35:12]
  assign _GEN_6076 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_6075); // @[FFT.scala 35:12]
  assign _GEN_6077 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_6076); // @[FFT.scala 35:12]
  assign _GEN_6078 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_6077); // @[FFT.scala 35:12]
  assign _GEN_6079 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_6078); // @[FFT.scala 35:12]
  assign _GEN_6130 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_6131 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_6130); // @[FFT.scala 34:12]
  assign _GEN_6132 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_6131); // @[FFT.scala 34:12]
  assign _GEN_6133 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_6132); // @[FFT.scala 34:12]
  assign _GEN_6134 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_6133); // @[FFT.scala 34:12]
  assign _GEN_6135 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_6134); // @[FFT.scala 34:12]
  assign _GEN_6138 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_6139 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_6138); // @[FFT.scala 35:12]
  assign _GEN_6140 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_6139); // @[FFT.scala 35:12]
  assign _GEN_6141 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_6140); // @[FFT.scala 35:12]
  assign _GEN_6142 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_6141); // @[FFT.scala 35:12]
  assign _GEN_6143 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_6142); // @[FFT.scala 35:12]
  assign _GEN_6170 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_6171 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_6170); // @[FFT.scala 34:12]
  assign _GEN_6174 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_6175 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_6174); // @[FFT.scala 35:12]
  assign io_dOut1_re = _T_3335_re; // @[FFT.scala 85:12]
  assign io_dOut1_im = _T_3335_im; // @[FFT.scala 85:12]
  assign io_dOut2_re = _T_3336_re; // @[FFT.scala 86:12]
  assign io_dOut2_im = _T_3336_im; // @[FFT.scala 86:12]
  assign io_dout_valid = cntD2 == 11'h7ff; // @[FFT.scala 88:19]
  assign BRAM_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_addr = cnt[9:0]; // @[FFT.scala 64:19]
  assign Butterfly_io_in1_re = _T_1204_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_1204_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = out2_0_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = out2_0_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = _T_176[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = _T_176[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_1718_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_1718_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cntD1[9]; // @[Butterfly.scala 113:17]
  assign BRAM_1_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_1_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_1_addr = cnt[8:0]; // @[FFT.scala 64:19]
  assign Butterfly_1_io_in1_re = _T_2239_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_2239_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = _T_1723[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = _T_1723[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_2497_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_2497_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cntD1[8]; // @[Butterfly.scala 113:17]
  assign BRAM_2_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_2_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_2_addr = cnt[7:0]; // @[FFT.scala 64:19]
  assign Butterfly_2_io_in1_re = _T_2762_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_2762_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = _T_2502[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = _T_2502[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_2892_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_2892_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cntD1[7]; // @[Butterfly.scala 113:17]
  assign BRAM_3_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_3_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_3_addr = cnt[6:0]; // @[FFT.scala 64:19]
  assign Butterfly_3_io_in1_re = _T_3029_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_3029_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = _T_2897[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = _T_2897[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_3095_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_3095_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cntD1[6]; // @[Butterfly.scala 113:17]
  assign BRAM_4_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_4_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_4_addr = cnt[5:0]; // @[FFT.scala 64:19]
  assign Butterfly_4_io_in1_re = _T_3168_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_3168_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = _T_3100[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = _T_3100[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_3202_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_3202_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cntD1[5]; // @[Butterfly.scala 113:17]
  assign BRAM_5_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_5_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_5_addr = cnt[4:0]; // @[FFT.scala 64:19]
  assign Butterfly_5_io_in1_re = _T_3243_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_3243_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = _T_3207[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = _T_3207[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_3261_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_3261_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cntD1[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_3282_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_3282_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_6063); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_6079); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_3292_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_3292_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cntD1[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_7_io_in1_re = _T_3305_re; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in1_im = _T_3305_im; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_6135); // @[Butterfly.scala 92:16]
  assign Butterfly_7_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_6143); // @[Butterfly.scala 92:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in2_re = _T_3311_re; // @[Butterfly.scala 112:17]
  assign Switch_7_io_in2_im = _T_3311_im; // @[Butterfly.scala 112:17]
  assign Switch_7_io_sel = cntD1[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_8_io_in1_re = _T_3320_re; // @[Butterfly.scala 90:17]
  assign Butterfly_8_io_in1_im = _T_3320_im; // @[Butterfly.scala 90:17]
  assign Butterfly_8_io_in2_re = Switch_7_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_8_io_in2_im = Switch_7_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_8_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_6171); // @[Butterfly.scala 92:16]
  assign Butterfly_8_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_6175); // @[Butterfly.scala 92:16]
  assign Switch_8_io_in1_re = Butterfly_8_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_8_io_in1_im = Butterfly_8_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_8_io_in2_re = _T_3324_re; // @[Butterfly.scala 112:17]
  assign Switch_8_io_in2_im = _T_3324_im; // @[Butterfly.scala 112:17]
  assign Switch_8_io_sel = cntD1[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_9_io_in1_re = _T_3331_re; // @[Butterfly.scala 90:17]
  assign Butterfly_9_io_in1_im = _T_3331_im; // @[Butterfly.scala 90:17]
  assign Butterfly_9_io_in2_re = Switch_8_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_9_io_in2_im = Switch_8_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_9_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_9_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_9_io_in1_re = Butterfly_9_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_9_io_in1_im = Butterfly_9_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_9_io_in2_re = _T_3334_re; // @[Butterfly.scala 112:17]
  assign Switch_9_io_in2_im = _T_3334_im; // @[Butterfly.scala 112:17]
  assign Switch_9_io_sel = cntD1[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_9_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_9_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_9_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_9_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntD1 = _RAND_1[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cntD2 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out1_0_re = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out1_0_im = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out2_0_re = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out2_0_im = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_181_re = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_181_im = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_182_re = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_182_im = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_183_re = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_183_im = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_184_re = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_184_im = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_185_re = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_185_im = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_186_re = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_186_im = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_187_re = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_187_im = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_188_re = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_188_im = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_189_re = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_189_im = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_190_re = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_190_im = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_191_re = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_191_im = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_192_re = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_192_im = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_193_re = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_193_im = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_194_re = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_194_im = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_195_re = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_195_im = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_196_re = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_196_im = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_197_re = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_197_im = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_198_re = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_198_im = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_199_re = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_199_im = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_200_re = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_200_im = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_201_re = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_201_im = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_202_re = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_202_im = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_203_re = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_203_im = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_204_re = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_204_im = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_205_re = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_205_im = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_206_re = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_206_im = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_207_re = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_207_im = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_208_re = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_208_im = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_209_re = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_209_im = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_210_re = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_210_im = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_211_re = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_211_im = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_212_re = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_212_im = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_213_re = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_213_im = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_214_re = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_214_im = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_215_re = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_215_im = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_216_re = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_216_im = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_217_re = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_217_im = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_218_re = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_218_im = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_219_re = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_219_im = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_220_re = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_220_im = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_221_re = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_221_im = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_222_re = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_222_im = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_223_re = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_223_im = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_224_re = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_224_im = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_225_re = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_225_im = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_226_re = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_226_im = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_227_re = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_227_im = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_228_re = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_228_im = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_229_re = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_229_im = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_230_re = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_230_im = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_231_re = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_231_im = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_232_re = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_232_im = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_233_re = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_233_im = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_234_re = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_234_im = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_235_re = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_235_im = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_236_re = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_236_im = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_237_re = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_237_im = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_238_re = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_238_im = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_239_re = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_239_im = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_240_re = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_240_im = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_241_re = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_241_im = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_242_re = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_242_im = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_243_re = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_243_im = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_244_re = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_244_im = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_245_re = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_245_im = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_246_re = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_246_im = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_247_re = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_247_im = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_248_re = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_248_im = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_249_re = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_249_im = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_250_re = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_250_im = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_251_re = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_251_im = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_252_re = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_252_im = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_253_re = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_253_im = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_254_re = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_254_im = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_255_re = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_255_im = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_256_re = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_256_im = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_257_re = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_257_im = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_258_re = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_258_im = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_259_re = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_259_im = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_260_re = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_260_im = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_261_re = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_261_im = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_262_re = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_262_im = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_263_re = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_263_im = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_264_re = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_264_im = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_265_re = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_265_im = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_266_re = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_266_im = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_267_re = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_267_im = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_268_re = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_268_im = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_269_re = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_269_im = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_270_re = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_270_im = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_271_re = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_271_im = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_272_re = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_272_im = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_273_re = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_273_im = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_274_re = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_274_im = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_275_re = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_275_im = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_276_re = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_276_im = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_277_re = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_277_im = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_278_re = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_278_im = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_279_re = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_279_im = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_280_re = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_280_im = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_281_re = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_281_im = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_282_re = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_282_im = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_283_re = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_283_im = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_284_re = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_284_im = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_285_re = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_285_im = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_286_re = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_286_im = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_287_re = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_287_im = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_288_re = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_288_im = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_289_re = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_289_im = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_290_re = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_290_im = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_291_re = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_291_im = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_292_re = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_292_im = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_293_re = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_293_im = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_294_re = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_294_im = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_295_re = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_295_im = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_296_re = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_296_im = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_297_re = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_297_im = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_298_re = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_298_im = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_299_re = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_299_im = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_300_re = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_300_im = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_301_re = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_301_im = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_302_re = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_302_im = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_303_re = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_303_im = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_304_re = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_304_im = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_305_re = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_305_im = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_306_re = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_306_im = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_307_re = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_307_im = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_308_re = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_308_im = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_309_re = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_309_im = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_310_re = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_310_im = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_311_re = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_311_im = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_312_re = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_312_im = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_313_re = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_313_im = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_314_re = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_314_im = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_315_re = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_315_im = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_316_re = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_316_im = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_317_re = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_317_im = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_318_re = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_318_im = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_319_re = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_319_im = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_320_re = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_320_im = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_321_re = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_321_im = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_322_re = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_322_im = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_323_re = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_323_im = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_324_re = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_324_im = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_325_re = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_325_im = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_326_re = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_326_im = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_327_re = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_327_im = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_328_re = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_328_im = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_329_re = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_329_im = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_330_re = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_330_im = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_331_re = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_331_im = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_332_re = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_332_im = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_333_re = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_333_im = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_334_re = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_334_im = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_335_re = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_335_im = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_336_re = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_336_im = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_337_re = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_337_im = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_338_re = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_338_im = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_339_re = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_339_im = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_340_re = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_340_im = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_341_re = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_341_im = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_342_re = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_342_im = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_343_re = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_343_im = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_344_re = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_344_im = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_345_re = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_345_im = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_346_re = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_346_im = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_347_re = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_347_im = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_348_re = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_348_im = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_349_re = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_349_im = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_350_re = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_350_im = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_351_re = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_351_im = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_352_re = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_352_im = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_353_re = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_353_im = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_354_re = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_354_im = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_355_re = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_355_im = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_356_re = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_356_im = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_357_re = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_357_im = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_358_re = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_358_im = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_359_re = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_359_im = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_360_re = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_360_im = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_361_re = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_361_im = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_362_re = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_362_im = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_363_re = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_363_im = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_364_re = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_364_im = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_365_re = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_365_im = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_366_re = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_366_im = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_367_re = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_367_im = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_368_re = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_368_im = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_369_re = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_369_im = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_370_re = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_370_im = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_371_re = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_371_im = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_372_re = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_372_im = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_373_re = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_373_im = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_374_re = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_374_im = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_375_re = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_375_im = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_376_re = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_376_im = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_377_re = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_377_im = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_378_re = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_378_im = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_379_re = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_379_im = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_380_re = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_380_im = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_381_re = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_381_im = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_382_re = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_382_im = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_383_re = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_383_im = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_384_re = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_384_im = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_385_re = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_385_im = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_386_re = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_386_im = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_387_re = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_387_im = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_388_re = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_388_im = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_389_re = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_389_im = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_390_re = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_390_im = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_391_re = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_391_im = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_392_re = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_392_im = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_393_re = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_393_im = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_394_re = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_394_im = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_395_re = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_395_im = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_396_re = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_396_im = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_397_re = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_397_im = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_398_re = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_398_im = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_399_re = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_399_im = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_400_re = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_400_im = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_401_re = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_401_im = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_402_re = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_402_im = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_403_re = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_403_im = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_404_re = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_404_im = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_405_re = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_405_im = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_406_re = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_406_im = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_407_re = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_407_im = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_408_re = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_408_im = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_409_re = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_409_im = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_410_re = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_410_im = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_411_re = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_411_im = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_412_re = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_412_im = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_413_re = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_413_im = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_414_re = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_414_im = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_415_re = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_415_im = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_416_re = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_416_im = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_417_re = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_417_im = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_418_re = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_418_im = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_419_re = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_419_im = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_420_re = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_420_im = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_421_re = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_421_im = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_422_re = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_422_im = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_423_re = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_423_im = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_424_re = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_424_im = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_425_re = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_425_im = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_426_re = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_426_im = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_427_re = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_427_im = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_428_re = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_428_im = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_429_re = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_429_im = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_430_re = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_430_im = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_431_re = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_431_im = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_432_re = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_432_im = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_433_re = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_433_im = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_434_re = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_434_im = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_435_re = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_435_im = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_436_re = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_436_im = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_437_re = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_437_im = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_438_re = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_438_im = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_439_re = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_439_im = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_440_re = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_440_im = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_441_re = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_441_im = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_442_re = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_442_im = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_443_re = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_443_im = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_444_re = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_444_im = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_445_re = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_445_im = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_446_re = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_446_im = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_447_re = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_447_im = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_448_re = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_448_im = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_449_re = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_449_im = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_450_re = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_450_im = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_451_re = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_451_im = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_452_re = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_452_im = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_453_re = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_453_im = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_454_re = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_454_im = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_455_re = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_455_im = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_456_re = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_456_im = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_457_re = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_457_im = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_458_re = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_458_im = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_459_re = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_459_im = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_460_re = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_460_im = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_461_re = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_461_im = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_462_re = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_462_im = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_463_re = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_463_im = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_464_re = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_464_im = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_465_re = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_465_im = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_466_re = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_466_im = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_467_re = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_467_im = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_468_re = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_468_im = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_469_re = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_469_im = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_470_re = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_470_im = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_471_re = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_471_im = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_472_re = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_472_im = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_473_re = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_473_im = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_474_re = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_474_im = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_475_re = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_475_im = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_476_re = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_476_im = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_477_re = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_477_im = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_478_re = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_478_im = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_479_re = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_479_im = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_480_re = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_480_im = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_481_re = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_481_im = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_482_re = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_482_im = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_483_re = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_483_im = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_484_re = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_484_im = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_485_re = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_485_im = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_486_re = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_486_im = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_487_re = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_487_im = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_488_re = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_488_im = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_489_re = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_489_im = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_490_re = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_490_im = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_491_re = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_491_im = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_492_re = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_492_im = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_493_re = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_493_im = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_494_re = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_494_im = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_495_re = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_495_im = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_496_re = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_496_im = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_497_re = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_497_im = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_498_re = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_498_im = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_499_re = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_499_im = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_500_re = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_500_im = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_501_re = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_501_im = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_502_re = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_502_im = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_503_re = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_503_im = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_504_re = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_504_im = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_505_re = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_505_im = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_506_re = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_506_im = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_507_re = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_507_im = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_508_re = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_508_im = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_509_re = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_509_im = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_510_re = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_510_im = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_511_re = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_511_im = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_512_re = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_512_im = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_513_re = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_513_im = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_514_re = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_514_im = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_515_re = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_515_im = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_516_re = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_516_im = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_517_re = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_517_im = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_518_re = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_518_im = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_519_re = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_519_im = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_520_re = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_520_im = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_521_re = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_521_im = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_522_re = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_522_im = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_523_re = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_523_im = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_524_re = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_524_im = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_525_re = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_525_im = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_526_re = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_526_im = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_527_re = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_527_im = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_528_re = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_528_im = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_529_re = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_529_im = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_530_re = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_530_im = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_531_re = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_531_im = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_532_re = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_532_im = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_533_re = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_533_im = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_534_re = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_534_im = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_535_re = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_535_im = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_536_re = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_536_im = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_537_re = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_537_im = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_538_re = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_538_im = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_539_re = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_539_im = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_540_re = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_540_im = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_541_re = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_541_im = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_542_re = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_542_im = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_543_re = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_543_im = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_544_re = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_544_im = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_545_re = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_545_im = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_546_re = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_546_im = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_547_re = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_547_im = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_548_re = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_548_im = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_549_re = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_549_im = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_550_re = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_550_im = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_551_re = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_551_im = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_552_re = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_552_im = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_553_re = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_553_im = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_554_re = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_554_im = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_555_re = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_555_im = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_556_re = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_556_im = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_557_re = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_557_im = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_558_re = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_558_im = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_559_re = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_559_im = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_560_re = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_560_im = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_561_re = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_561_im = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_562_re = _RAND_769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_562_im = _RAND_770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_563_re = _RAND_771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_563_im = _RAND_772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_564_re = _RAND_773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_564_im = _RAND_774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_565_re = _RAND_775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_565_im = _RAND_776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_566_re = _RAND_777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_566_im = _RAND_778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_567_re = _RAND_779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_567_im = _RAND_780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_568_re = _RAND_781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_568_im = _RAND_782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_569_re = _RAND_783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_569_im = _RAND_784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_570_re = _RAND_785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_570_im = _RAND_786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_571_re = _RAND_787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_571_im = _RAND_788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_572_re = _RAND_789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_572_im = _RAND_790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_573_re = _RAND_791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_573_im = _RAND_792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_574_re = _RAND_793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_574_im = _RAND_794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_575_re = _RAND_795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_575_im = _RAND_796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_576_re = _RAND_797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_576_im = _RAND_798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_577_re = _RAND_799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_577_im = _RAND_800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_578_re = _RAND_801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_578_im = _RAND_802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_579_re = _RAND_803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_579_im = _RAND_804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_580_re = _RAND_805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_580_im = _RAND_806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_581_re = _RAND_807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_581_im = _RAND_808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_582_re = _RAND_809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_582_im = _RAND_810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_583_re = _RAND_811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_583_im = _RAND_812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_584_re = _RAND_813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_584_im = _RAND_814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_585_re = _RAND_815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_585_im = _RAND_816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_586_re = _RAND_817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_586_im = _RAND_818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_587_re = _RAND_819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_587_im = _RAND_820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_588_re = _RAND_821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_588_im = _RAND_822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_589_re = _RAND_823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_589_im = _RAND_824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_590_re = _RAND_825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_590_im = _RAND_826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_591_re = _RAND_827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_591_im = _RAND_828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_592_re = _RAND_829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_592_im = _RAND_830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_593_re = _RAND_831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_593_im = _RAND_832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_594_re = _RAND_833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_594_im = _RAND_834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_595_re = _RAND_835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_595_im = _RAND_836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_596_re = _RAND_837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_596_im = _RAND_838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_597_re = _RAND_839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_597_im = _RAND_840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_598_re = _RAND_841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_598_im = _RAND_842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_599_re = _RAND_843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_599_im = _RAND_844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_600_re = _RAND_845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_600_im = _RAND_846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_601_re = _RAND_847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_601_im = _RAND_848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_602_re = _RAND_849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_602_im = _RAND_850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_603_re = _RAND_851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_603_im = _RAND_852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_604_re = _RAND_853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_604_im = _RAND_854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_605_re = _RAND_855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_605_im = _RAND_856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_606_re = _RAND_857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_606_im = _RAND_858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_607_re = _RAND_859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_607_im = _RAND_860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_608_re = _RAND_861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_608_im = _RAND_862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_609_re = _RAND_863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_609_im = _RAND_864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_610_re = _RAND_865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_610_im = _RAND_866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_611_re = _RAND_867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_611_im = _RAND_868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_612_re = _RAND_869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_612_im = _RAND_870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_613_re = _RAND_871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_613_im = _RAND_872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_614_re = _RAND_873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_614_im = _RAND_874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_615_re = _RAND_875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_615_im = _RAND_876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_616_re = _RAND_877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_616_im = _RAND_878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_617_re = _RAND_879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_617_im = _RAND_880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_618_re = _RAND_881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_618_im = _RAND_882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_619_re = _RAND_883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_619_im = _RAND_884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_620_re = _RAND_885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_620_im = _RAND_886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_621_re = _RAND_887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_621_im = _RAND_888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_622_re = _RAND_889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_622_im = _RAND_890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_623_re = _RAND_891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_623_im = _RAND_892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_624_re = _RAND_893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_624_im = _RAND_894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_625_re = _RAND_895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_625_im = _RAND_896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_626_re = _RAND_897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_626_im = _RAND_898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_627_re = _RAND_899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_627_im = _RAND_900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_628_re = _RAND_901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_628_im = _RAND_902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_629_re = _RAND_903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_629_im = _RAND_904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_630_re = _RAND_905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_630_im = _RAND_906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_631_re = _RAND_907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_631_im = _RAND_908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_632_re = _RAND_909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_632_im = _RAND_910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_633_re = _RAND_911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_633_im = _RAND_912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_634_re = _RAND_913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_634_im = _RAND_914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_635_re = _RAND_915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_635_im = _RAND_916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_636_re = _RAND_917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_636_im = _RAND_918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_637_re = _RAND_919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_637_im = _RAND_920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_638_re = _RAND_921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_638_im = _RAND_922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_639_re = _RAND_923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_639_im = _RAND_924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_640_re = _RAND_925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_640_im = _RAND_926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_641_re = _RAND_927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_641_im = _RAND_928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_642_re = _RAND_929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_642_im = _RAND_930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_643_re = _RAND_931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_643_im = _RAND_932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_644_re = _RAND_933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_644_im = _RAND_934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_645_re = _RAND_935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_645_im = _RAND_936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_646_re = _RAND_937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_646_im = _RAND_938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_647_re = _RAND_939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_647_im = _RAND_940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_648_re = _RAND_941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_648_im = _RAND_942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_649_re = _RAND_943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_649_im = _RAND_944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_650_re = _RAND_945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_650_im = _RAND_946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_651_re = _RAND_947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_651_im = _RAND_948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_652_re = _RAND_949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_652_im = _RAND_950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_653_re = _RAND_951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_653_im = _RAND_952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_654_re = _RAND_953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_654_im = _RAND_954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_655_re = _RAND_955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_655_im = _RAND_956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_656_re = _RAND_957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_656_im = _RAND_958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_657_re = _RAND_959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_657_im = _RAND_960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_658_re = _RAND_961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_658_im = _RAND_962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_659_re = _RAND_963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_659_im = _RAND_964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_660_re = _RAND_965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_660_im = _RAND_966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_661_re = _RAND_967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_661_im = _RAND_968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_662_re = _RAND_969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_662_im = _RAND_970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_663_re = _RAND_971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_663_im = _RAND_972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_664_re = _RAND_973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_664_im = _RAND_974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_665_re = _RAND_975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_665_im = _RAND_976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_666_re = _RAND_977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_666_im = _RAND_978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_667_re = _RAND_979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_667_im = _RAND_980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_668_re = _RAND_981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_668_im = _RAND_982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_669_re = _RAND_983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_669_im = _RAND_984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_670_re = _RAND_985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_670_im = _RAND_986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_671_re = _RAND_987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_671_im = _RAND_988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_672_re = _RAND_989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_672_im = _RAND_990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_673_re = _RAND_991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_673_im = _RAND_992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_674_re = _RAND_993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_674_im = _RAND_994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_675_re = _RAND_995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_675_im = _RAND_996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_676_re = _RAND_997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_676_im = _RAND_998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_677_re = _RAND_999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_677_im = _RAND_1000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_678_re = _RAND_1001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_678_im = _RAND_1002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_679_re = _RAND_1003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_679_im = _RAND_1004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_680_re = _RAND_1005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_680_im = _RAND_1006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_681_re = _RAND_1007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_681_im = _RAND_1008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_682_re = _RAND_1009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_682_im = _RAND_1010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_683_re = _RAND_1011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_683_im = _RAND_1012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_684_re = _RAND_1013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_684_im = _RAND_1014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_685_re = _RAND_1015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_685_im = _RAND_1016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_686_re = _RAND_1017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_686_im = _RAND_1018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_687_re = _RAND_1019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_687_im = _RAND_1020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_688_re = _RAND_1021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_688_im = _RAND_1022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_689_re = _RAND_1023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_689_im = _RAND_1024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_690_re = _RAND_1025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_690_im = _RAND_1026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_691_re = _RAND_1027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_691_im = _RAND_1028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_692_re = _RAND_1029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_692_im = _RAND_1030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_693_re = _RAND_1031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_693_im = _RAND_1032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_694_re = _RAND_1033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_694_im = _RAND_1034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_695_re = _RAND_1035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_695_im = _RAND_1036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_696_re = _RAND_1037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_696_im = _RAND_1038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_697_re = _RAND_1039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_697_im = _RAND_1040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_698_re = _RAND_1041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_698_im = _RAND_1042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_699_re = _RAND_1043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_699_im = _RAND_1044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_700_re = _RAND_1045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_700_im = _RAND_1046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_701_re = _RAND_1047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_701_im = _RAND_1048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_702_re = _RAND_1049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_702_im = _RAND_1050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_703_re = _RAND_1051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_703_im = _RAND_1052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_704_re = _RAND_1053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_704_im = _RAND_1054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_705_re = _RAND_1055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_705_im = _RAND_1056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_706_re = _RAND_1057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_706_im = _RAND_1058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_707_re = _RAND_1059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_707_im = _RAND_1060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_708_re = _RAND_1061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_708_im = _RAND_1062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_709_re = _RAND_1063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_709_im = _RAND_1064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_710_re = _RAND_1065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_710_im = _RAND_1066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_711_re = _RAND_1067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_711_im = _RAND_1068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_712_re = _RAND_1069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_712_im = _RAND_1070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_713_re = _RAND_1071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_713_im = _RAND_1072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_714_re = _RAND_1073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_714_im = _RAND_1074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_715_re = _RAND_1075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_715_im = _RAND_1076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_716_re = _RAND_1077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_716_im = _RAND_1078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_717_re = _RAND_1079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_717_im = _RAND_1080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_718_re = _RAND_1081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_718_im = _RAND_1082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_719_re = _RAND_1083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_719_im = _RAND_1084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_720_re = _RAND_1085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_720_im = _RAND_1086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_721_re = _RAND_1087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_721_im = _RAND_1088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_722_re = _RAND_1089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_722_im = _RAND_1090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_723_re = _RAND_1091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_723_im = _RAND_1092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_724_re = _RAND_1093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_724_im = _RAND_1094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_725_re = _RAND_1095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_725_im = _RAND_1096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_726_re = _RAND_1097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_726_im = _RAND_1098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_727_re = _RAND_1099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_727_im = _RAND_1100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_728_re = _RAND_1101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_728_im = _RAND_1102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_729_re = _RAND_1103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_729_im = _RAND_1104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_730_re = _RAND_1105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_730_im = _RAND_1106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_731_re = _RAND_1107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_731_im = _RAND_1108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_732_re = _RAND_1109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_732_im = _RAND_1110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_733_re = _RAND_1111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_733_im = _RAND_1112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_734_re = _RAND_1113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_734_im = _RAND_1114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_735_re = _RAND_1115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_735_im = _RAND_1116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_736_re = _RAND_1117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_736_im = _RAND_1118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_737_re = _RAND_1119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_737_im = _RAND_1120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_738_re = _RAND_1121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_738_im = _RAND_1122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_739_re = _RAND_1123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_739_im = _RAND_1124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_740_re = _RAND_1125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_740_im = _RAND_1126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_741_re = _RAND_1127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_741_im = _RAND_1128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_742_re = _RAND_1129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_742_im = _RAND_1130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_743_re = _RAND_1131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_743_im = _RAND_1132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_744_re = _RAND_1133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_744_im = _RAND_1134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_745_re = _RAND_1135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_745_im = _RAND_1136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_746_re = _RAND_1137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_746_im = _RAND_1138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_747_re = _RAND_1139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_747_im = _RAND_1140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_748_re = _RAND_1141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_748_im = _RAND_1142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_749_re = _RAND_1143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_749_im = _RAND_1144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_750_re = _RAND_1145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_750_im = _RAND_1146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_751_re = _RAND_1147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_751_im = _RAND_1148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_752_re = _RAND_1149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_752_im = _RAND_1150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_753_re = _RAND_1151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_753_im = _RAND_1152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_754_re = _RAND_1153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_754_im = _RAND_1154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_755_re = _RAND_1155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_755_im = _RAND_1156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_756_re = _RAND_1157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_756_im = _RAND_1158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_757_re = _RAND_1159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_757_im = _RAND_1160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_758_re = _RAND_1161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_758_im = _RAND_1162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_759_re = _RAND_1163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_759_im = _RAND_1164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_760_re = _RAND_1165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_760_im = _RAND_1166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_761_re = _RAND_1167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_761_im = _RAND_1168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_762_re = _RAND_1169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_762_im = _RAND_1170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_763_re = _RAND_1171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_763_im = _RAND_1172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_764_re = _RAND_1173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_764_im = _RAND_1174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_765_re = _RAND_1175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_765_im = _RAND_1176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_766_re = _RAND_1177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_766_im = _RAND_1178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_767_re = _RAND_1179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_767_im = _RAND_1180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_768_re = _RAND_1181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_768_im = _RAND_1182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_769_re = _RAND_1183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_769_im = _RAND_1184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_770_re = _RAND_1185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_770_im = _RAND_1186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_771_re = _RAND_1187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_771_im = _RAND_1188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_772_re = _RAND_1189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_772_im = _RAND_1190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_773_re = _RAND_1191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_773_im = _RAND_1192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_774_re = _RAND_1193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_774_im = _RAND_1194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_775_re = _RAND_1195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_775_im = _RAND_1196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_776_re = _RAND_1197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_776_im = _RAND_1198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_777_re = _RAND_1199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_777_im = _RAND_1200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_778_re = _RAND_1201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_778_im = _RAND_1202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_779_re = _RAND_1203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_779_im = _RAND_1204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_780_re = _RAND_1205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_780_im = _RAND_1206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_781_re = _RAND_1207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_781_im = _RAND_1208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_782_re = _RAND_1209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_782_im = _RAND_1210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_783_re = _RAND_1211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_783_im = _RAND_1212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_784_re = _RAND_1213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_784_im = _RAND_1214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_785_re = _RAND_1215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_785_im = _RAND_1216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_786_re = _RAND_1217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_786_im = _RAND_1218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_787_re = _RAND_1219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_787_im = _RAND_1220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_788_re = _RAND_1221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_788_im = _RAND_1222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_789_re = _RAND_1223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_789_im = _RAND_1224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_790_re = _RAND_1225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_790_im = _RAND_1226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_791_re = _RAND_1227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_791_im = _RAND_1228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_792_re = _RAND_1229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_792_im = _RAND_1230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_793_re = _RAND_1231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_793_im = _RAND_1232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_794_re = _RAND_1233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_794_im = _RAND_1234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_795_re = _RAND_1235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_795_im = _RAND_1236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_796_re = _RAND_1237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_796_im = _RAND_1238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_797_re = _RAND_1239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_797_im = _RAND_1240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_798_re = _RAND_1241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_798_im = _RAND_1242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_799_re = _RAND_1243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_799_im = _RAND_1244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_800_re = _RAND_1245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_800_im = _RAND_1246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_801_re = _RAND_1247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_801_im = _RAND_1248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_802_re = _RAND_1249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_802_im = _RAND_1250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_803_re = _RAND_1251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  _T_803_im = _RAND_1252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  _T_804_re = _RAND_1253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  _T_804_im = _RAND_1254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  _T_805_re = _RAND_1255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  _T_805_im = _RAND_1256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  _T_806_re = _RAND_1257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  _T_806_im = _RAND_1258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  _T_807_re = _RAND_1259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  _T_807_im = _RAND_1260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  _T_808_re = _RAND_1261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  _T_808_im = _RAND_1262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  _T_809_re = _RAND_1263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  _T_809_im = _RAND_1264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  _T_810_re = _RAND_1265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  _T_810_im = _RAND_1266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  _T_811_re = _RAND_1267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  _T_811_im = _RAND_1268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  _T_812_re = _RAND_1269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  _T_812_im = _RAND_1270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  _T_813_re = _RAND_1271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  _T_813_im = _RAND_1272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  _T_814_re = _RAND_1273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  _T_814_im = _RAND_1274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  _T_815_re = _RAND_1275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  _T_815_im = _RAND_1276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  _T_816_re = _RAND_1277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  _T_816_im = _RAND_1278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  _T_817_re = _RAND_1279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  _T_817_im = _RAND_1280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  _T_818_re = _RAND_1281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  _T_818_im = _RAND_1282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  _T_819_re = _RAND_1283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  _T_819_im = _RAND_1284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  _T_820_re = _RAND_1285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  _T_820_im = _RAND_1286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  _T_821_re = _RAND_1287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  _T_821_im = _RAND_1288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  _T_822_re = _RAND_1289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  _T_822_im = _RAND_1290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  _T_823_re = _RAND_1291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  _T_823_im = _RAND_1292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  _T_824_re = _RAND_1293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  _T_824_im = _RAND_1294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  _T_825_re = _RAND_1295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  _T_825_im = _RAND_1296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  _T_826_re = _RAND_1297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  _T_826_im = _RAND_1298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  _T_827_re = _RAND_1299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  _T_827_im = _RAND_1300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  _T_828_re = _RAND_1301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  _T_828_im = _RAND_1302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  _T_829_re = _RAND_1303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  _T_829_im = _RAND_1304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  _T_830_re = _RAND_1305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  _T_830_im = _RAND_1306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  _T_831_re = _RAND_1307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  _T_831_im = _RAND_1308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  _T_832_re = _RAND_1309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  _T_832_im = _RAND_1310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  _T_833_re = _RAND_1311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  _T_833_im = _RAND_1312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  _T_834_re = _RAND_1313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  _T_834_im = _RAND_1314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  _T_835_re = _RAND_1315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  _T_835_im = _RAND_1316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  _T_836_re = _RAND_1317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  _T_836_im = _RAND_1318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  _T_837_re = _RAND_1319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  _T_837_im = _RAND_1320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  _T_838_re = _RAND_1321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  _T_838_im = _RAND_1322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  _T_839_re = _RAND_1323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  _T_839_im = _RAND_1324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  _T_840_re = _RAND_1325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  _T_840_im = _RAND_1326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  _T_841_re = _RAND_1327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  _T_841_im = _RAND_1328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  _T_842_re = _RAND_1329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  _T_842_im = _RAND_1330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  _T_843_re = _RAND_1331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  _T_843_im = _RAND_1332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  _T_844_re = _RAND_1333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  _T_844_im = _RAND_1334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  _T_845_re = _RAND_1335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  _T_845_im = _RAND_1336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  _T_846_re = _RAND_1337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  _T_846_im = _RAND_1338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  _T_847_re = _RAND_1339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  _T_847_im = _RAND_1340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  _T_848_re = _RAND_1341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  _T_848_im = _RAND_1342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  _T_849_re = _RAND_1343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  _T_849_im = _RAND_1344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  _T_850_re = _RAND_1345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  _T_850_im = _RAND_1346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  _T_851_re = _RAND_1347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  _T_851_im = _RAND_1348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  _T_852_re = _RAND_1349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  _T_852_im = _RAND_1350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  _T_853_re = _RAND_1351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  _T_853_im = _RAND_1352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  _T_854_re = _RAND_1353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  _T_854_im = _RAND_1354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  _T_855_re = _RAND_1355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  _T_855_im = _RAND_1356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  _T_856_re = _RAND_1357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  _T_856_im = _RAND_1358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  _T_857_re = _RAND_1359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  _T_857_im = _RAND_1360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  _T_858_re = _RAND_1361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  _T_858_im = _RAND_1362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  _T_859_re = _RAND_1363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  _T_859_im = _RAND_1364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  _T_860_re = _RAND_1365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  _T_860_im = _RAND_1366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  _T_861_re = _RAND_1367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  _T_861_im = _RAND_1368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  _T_862_re = _RAND_1369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  _T_862_im = _RAND_1370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  _T_863_re = _RAND_1371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  _T_863_im = _RAND_1372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  _T_864_re = _RAND_1373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  _T_864_im = _RAND_1374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  _T_865_re = _RAND_1375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  _T_865_im = _RAND_1376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  _T_866_re = _RAND_1377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  _T_866_im = _RAND_1378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  _T_867_re = _RAND_1379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  _T_867_im = _RAND_1380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  _T_868_re = _RAND_1381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  _T_868_im = _RAND_1382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  _T_869_re = _RAND_1383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  _T_869_im = _RAND_1384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  _T_870_re = _RAND_1385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  _T_870_im = _RAND_1386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  _T_871_re = _RAND_1387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  _T_871_im = _RAND_1388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  _T_872_re = _RAND_1389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  _T_872_im = _RAND_1390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  _T_873_re = _RAND_1391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  _T_873_im = _RAND_1392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  _T_874_re = _RAND_1393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  _T_874_im = _RAND_1394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  _T_875_re = _RAND_1395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  _T_875_im = _RAND_1396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  _T_876_re = _RAND_1397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  _T_876_im = _RAND_1398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  _T_877_re = _RAND_1399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  _T_877_im = _RAND_1400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  _T_878_re = _RAND_1401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  _T_878_im = _RAND_1402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  _T_879_re = _RAND_1403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  _T_879_im = _RAND_1404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  _T_880_re = _RAND_1405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  _T_880_im = _RAND_1406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  _T_881_re = _RAND_1407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  _T_881_im = _RAND_1408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  _T_882_re = _RAND_1409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  _T_882_im = _RAND_1410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  _T_883_re = _RAND_1411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  _T_883_im = _RAND_1412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  _T_884_re = _RAND_1413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  _T_884_im = _RAND_1414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  _T_885_re = _RAND_1415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  _T_885_im = _RAND_1416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  _T_886_re = _RAND_1417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  _T_886_im = _RAND_1418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  _T_887_re = _RAND_1419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  _T_887_im = _RAND_1420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  _T_888_re = _RAND_1421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  _T_888_im = _RAND_1422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  _T_889_re = _RAND_1423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  _T_889_im = _RAND_1424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  _T_890_re = _RAND_1425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  _T_890_im = _RAND_1426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  _T_891_re = _RAND_1427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  _T_891_im = _RAND_1428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  _T_892_re = _RAND_1429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  _T_892_im = _RAND_1430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  _T_893_re = _RAND_1431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  _T_893_im = _RAND_1432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  _T_894_re = _RAND_1433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  _T_894_im = _RAND_1434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  _T_895_re = _RAND_1435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  _T_895_im = _RAND_1436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  _T_896_re = _RAND_1437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  _T_896_im = _RAND_1438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  _T_897_re = _RAND_1439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  _T_897_im = _RAND_1440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  _T_898_re = _RAND_1441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  _T_898_im = _RAND_1442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  _T_899_re = _RAND_1443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  _T_899_im = _RAND_1444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  _T_900_re = _RAND_1445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  _T_900_im = _RAND_1446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  _T_901_re = _RAND_1447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  _T_901_im = _RAND_1448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  _T_902_re = _RAND_1449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  _T_902_im = _RAND_1450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  _T_903_re = _RAND_1451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  _T_903_im = _RAND_1452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  _T_904_re = _RAND_1453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  _T_904_im = _RAND_1454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  _T_905_re = _RAND_1455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  _T_905_im = _RAND_1456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  _T_906_re = _RAND_1457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  _T_906_im = _RAND_1458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  _T_907_re = _RAND_1459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  _T_907_im = _RAND_1460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  _T_908_re = _RAND_1461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  _T_908_im = _RAND_1462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  _T_909_re = _RAND_1463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  _T_909_im = _RAND_1464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  _T_910_re = _RAND_1465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  _T_910_im = _RAND_1466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  _T_911_re = _RAND_1467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  _T_911_im = _RAND_1468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  _T_912_re = _RAND_1469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  _T_912_im = _RAND_1470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  _T_913_re = _RAND_1471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  _T_913_im = _RAND_1472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  _T_914_re = _RAND_1473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  _T_914_im = _RAND_1474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  _T_915_re = _RAND_1475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  _T_915_im = _RAND_1476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  _T_916_re = _RAND_1477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  _T_916_im = _RAND_1478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  _T_917_re = _RAND_1479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  _T_917_im = _RAND_1480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  _T_918_re = _RAND_1481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  _T_918_im = _RAND_1482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  _T_919_re = _RAND_1483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  _T_919_im = _RAND_1484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  _T_920_re = _RAND_1485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  _T_920_im = _RAND_1486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  _T_921_re = _RAND_1487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  _T_921_im = _RAND_1488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  _T_922_re = _RAND_1489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  _T_922_im = _RAND_1490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  _T_923_re = _RAND_1491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  _T_923_im = _RAND_1492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  _T_924_re = _RAND_1493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  _T_924_im = _RAND_1494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  _T_925_re = _RAND_1495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  _T_925_im = _RAND_1496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  _T_926_re = _RAND_1497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  _T_926_im = _RAND_1498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  _T_927_re = _RAND_1499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  _T_927_im = _RAND_1500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  _T_928_re = _RAND_1501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  _T_928_im = _RAND_1502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  _T_929_re = _RAND_1503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  _T_929_im = _RAND_1504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  _T_930_re = _RAND_1505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  _T_930_im = _RAND_1506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  _T_931_re = _RAND_1507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  _T_931_im = _RAND_1508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  _T_932_re = _RAND_1509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  _T_932_im = _RAND_1510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  _T_933_re = _RAND_1511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  _T_933_im = _RAND_1512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  _T_934_re = _RAND_1513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  _T_934_im = _RAND_1514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  _T_935_re = _RAND_1515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  _T_935_im = _RAND_1516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  _T_936_re = _RAND_1517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  _T_936_im = _RAND_1518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  _T_937_re = _RAND_1519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  _T_937_im = _RAND_1520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  _T_938_re = _RAND_1521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  _T_938_im = _RAND_1522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  _T_939_re = _RAND_1523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  _T_939_im = _RAND_1524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  _T_940_re = _RAND_1525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  _T_940_im = _RAND_1526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  _T_941_re = _RAND_1527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  _T_941_im = _RAND_1528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  _T_942_re = _RAND_1529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  _T_942_im = _RAND_1530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  _T_943_re = _RAND_1531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  _T_943_im = _RAND_1532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  _T_944_re = _RAND_1533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  _T_944_im = _RAND_1534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  _T_945_re = _RAND_1535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  _T_945_im = _RAND_1536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  _T_946_re = _RAND_1537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  _T_946_im = _RAND_1538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  _T_947_re = _RAND_1539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  _T_947_im = _RAND_1540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  _T_948_re = _RAND_1541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  _T_948_im = _RAND_1542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1543 = {1{`RANDOM}};
  _T_949_re = _RAND_1543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1544 = {1{`RANDOM}};
  _T_949_im = _RAND_1544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1545 = {1{`RANDOM}};
  _T_950_re = _RAND_1545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1546 = {1{`RANDOM}};
  _T_950_im = _RAND_1546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1547 = {1{`RANDOM}};
  _T_951_re = _RAND_1547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1548 = {1{`RANDOM}};
  _T_951_im = _RAND_1548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1549 = {1{`RANDOM}};
  _T_952_re = _RAND_1549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1550 = {1{`RANDOM}};
  _T_952_im = _RAND_1550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1551 = {1{`RANDOM}};
  _T_953_re = _RAND_1551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1552 = {1{`RANDOM}};
  _T_953_im = _RAND_1552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1553 = {1{`RANDOM}};
  _T_954_re = _RAND_1553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1554 = {1{`RANDOM}};
  _T_954_im = _RAND_1554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1555 = {1{`RANDOM}};
  _T_955_re = _RAND_1555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1556 = {1{`RANDOM}};
  _T_955_im = _RAND_1556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1557 = {1{`RANDOM}};
  _T_956_re = _RAND_1557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1558 = {1{`RANDOM}};
  _T_956_im = _RAND_1558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1559 = {1{`RANDOM}};
  _T_957_re = _RAND_1559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1560 = {1{`RANDOM}};
  _T_957_im = _RAND_1560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1561 = {1{`RANDOM}};
  _T_958_re = _RAND_1561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1562 = {1{`RANDOM}};
  _T_958_im = _RAND_1562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1563 = {1{`RANDOM}};
  _T_959_re = _RAND_1563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1564 = {1{`RANDOM}};
  _T_959_im = _RAND_1564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1565 = {1{`RANDOM}};
  _T_960_re = _RAND_1565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1566 = {1{`RANDOM}};
  _T_960_im = _RAND_1566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1567 = {1{`RANDOM}};
  _T_961_re = _RAND_1567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1568 = {1{`RANDOM}};
  _T_961_im = _RAND_1568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1569 = {1{`RANDOM}};
  _T_962_re = _RAND_1569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1570 = {1{`RANDOM}};
  _T_962_im = _RAND_1570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1571 = {1{`RANDOM}};
  _T_963_re = _RAND_1571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1572 = {1{`RANDOM}};
  _T_963_im = _RAND_1572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1573 = {1{`RANDOM}};
  _T_964_re = _RAND_1573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1574 = {1{`RANDOM}};
  _T_964_im = _RAND_1574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1575 = {1{`RANDOM}};
  _T_965_re = _RAND_1575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1576 = {1{`RANDOM}};
  _T_965_im = _RAND_1576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1577 = {1{`RANDOM}};
  _T_966_re = _RAND_1577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1578 = {1{`RANDOM}};
  _T_966_im = _RAND_1578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1579 = {1{`RANDOM}};
  _T_967_re = _RAND_1579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1580 = {1{`RANDOM}};
  _T_967_im = _RAND_1580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1581 = {1{`RANDOM}};
  _T_968_re = _RAND_1581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1582 = {1{`RANDOM}};
  _T_968_im = _RAND_1582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1583 = {1{`RANDOM}};
  _T_969_re = _RAND_1583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1584 = {1{`RANDOM}};
  _T_969_im = _RAND_1584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1585 = {1{`RANDOM}};
  _T_970_re = _RAND_1585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1586 = {1{`RANDOM}};
  _T_970_im = _RAND_1586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1587 = {1{`RANDOM}};
  _T_971_re = _RAND_1587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1588 = {1{`RANDOM}};
  _T_971_im = _RAND_1588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1589 = {1{`RANDOM}};
  _T_972_re = _RAND_1589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1590 = {1{`RANDOM}};
  _T_972_im = _RAND_1590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1591 = {1{`RANDOM}};
  _T_973_re = _RAND_1591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1592 = {1{`RANDOM}};
  _T_973_im = _RAND_1592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1593 = {1{`RANDOM}};
  _T_974_re = _RAND_1593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1594 = {1{`RANDOM}};
  _T_974_im = _RAND_1594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1595 = {1{`RANDOM}};
  _T_975_re = _RAND_1595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1596 = {1{`RANDOM}};
  _T_975_im = _RAND_1596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1597 = {1{`RANDOM}};
  _T_976_re = _RAND_1597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1598 = {1{`RANDOM}};
  _T_976_im = _RAND_1598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1599 = {1{`RANDOM}};
  _T_977_re = _RAND_1599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1600 = {1{`RANDOM}};
  _T_977_im = _RAND_1600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1601 = {1{`RANDOM}};
  _T_978_re = _RAND_1601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1602 = {1{`RANDOM}};
  _T_978_im = _RAND_1602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1603 = {1{`RANDOM}};
  _T_979_re = _RAND_1603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1604 = {1{`RANDOM}};
  _T_979_im = _RAND_1604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1605 = {1{`RANDOM}};
  _T_980_re = _RAND_1605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1606 = {1{`RANDOM}};
  _T_980_im = _RAND_1606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1607 = {1{`RANDOM}};
  _T_981_re = _RAND_1607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1608 = {1{`RANDOM}};
  _T_981_im = _RAND_1608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1609 = {1{`RANDOM}};
  _T_982_re = _RAND_1609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1610 = {1{`RANDOM}};
  _T_982_im = _RAND_1610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1611 = {1{`RANDOM}};
  _T_983_re = _RAND_1611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1612 = {1{`RANDOM}};
  _T_983_im = _RAND_1612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1613 = {1{`RANDOM}};
  _T_984_re = _RAND_1613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1614 = {1{`RANDOM}};
  _T_984_im = _RAND_1614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1615 = {1{`RANDOM}};
  _T_985_re = _RAND_1615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1616 = {1{`RANDOM}};
  _T_985_im = _RAND_1616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1617 = {1{`RANDOM}};
  _T_986_re = _RAND_1617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1618 = {1{`RANDOM}};
  _T_986_im = _RAND_1618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1619 = {1{`RANDOM}};
  _T_987_re = _RAND_1619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1620 = {1{`RANDOM}};
  _T_987_im = _RAND_1620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1621 = {1{`RANDOM}};
  _T_988_re = _RAND_1621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1622 = {1{`RANDOM}};
  _T_988_im = _RAND_1622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1623 = {1{`RANDOM}};
  _T_989_re = _RAND_1623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1624 = {1{`RANDOM}};
  _T_989_im = _RAND_1624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1625 = {1{`RANDOM}};
  _T_990_re = _RAND_1625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1626 = {1{`RANDOM}};
  _T_990_im = _RAND_1626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1627 = {1{`RANDOM}};
  _T_991_re = _RAND_1627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1628 = {1{`RANDOM}};
  _T_991_im = _RAND_1628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1629 = {1{`RANDOM}};
  _T_992_re = _RAND_1629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1630 = {1{`RANDOM}};
  _T_992_im = _RAND_1630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1631 = {1{`RANDOM}};
  _T_993_re = _RAND_1631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1632 = {1{`RANDOM}};
  _T_993_im = _RAND_1632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1633 = {1{`RANDOM}};
  _T_994_re = _RAND_1633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1634 = {1{`RANDOM}};
  _T_994_im = _RAND_1634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1635 = {1{`RANDOM}};
  _T_995_re = _RAND_1635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1636 = {1{`RANDOM}};
  _T_995_im = _RAND_1636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1637 = {1{`RANDOM}};
  _T_996_re = _RAND_1637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1638 = {1{`RANDOM}};
  _T_996_im = _RAND_1638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1639 = {1{`RANDOM}};
  _T_997_re = _RAND_1639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1640 = {1{`RANDOM}};
  _T_997_im = _RAND_1640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1641 = {1{`RANDOM}};
  _T_998_re = _RAND_1641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1642 = {1{`RANDOM}};
  _T_998_im = _RAND_1642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1643 = {1{`RANDOM}};
  _T_999_re = _RAND_1643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1644 = {1{`RANDOM}};
  _T_999_im = _RAND_1644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1645 = {1{`RANDOM}};
  _T_1000_re = _RAND_1645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1646 = {1{`RANDOM}};
  _T_1000_im = _RAND_1646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1647 = {1{`RANDOM}};
  _T_1001_re = _RAND_1647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1648 = {1{`RANDOM}};
  _T_1001_im = _RAND_1648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1649 = {1{`RANDOM}};
  _T_1002_re = _RAND_1649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1650 = {1{`RANDOM}};
  _T_1002_im = _RAND_1650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1651 = {1{`RANDOM}};
  _T_1003_re = _RAND_1651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1652 = {1{`RANDOM}};
  _T_1003_im = _RAND_1652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1653 = {1{`RANDOM}};
  _T_1004_re = _RAND_1653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1654 = {1{`RANDOM}};
  _T_1004_im = _RAND_1654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1655 = {1{`RANDOM}};
  _T_1005_re = _RAND_1655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1656 = {1{`RANDOM}};
  _T_1005_im = _RAND_1656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1657 = {1{`RANDOM}};
  _T_1006_re = _RAND_1657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1658 = {1{`RANDOM}};
  _T_1006_im = _RAND_1658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1659 = {1{`RANDOM}};
  _T_1007_re = _RAND_1659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1660 = {1{`RANDOM}};
  _T_1007_im = _RAND_1660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1661 = {1{`RANDOM}};
  _T_1008_re = _RAND_1661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1662 = {1{`RANDOM}};
  _T_1008_im = _RAND_1662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1663 = {1{`RANDOM}};
  _T_1009_re = _RAND_1663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1664 = {1{`RANDOM}};
  _T_1009_im = _RAND_1664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1665 = {1{`RANDOM}};
  _T_1010_re = _RAND_1665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1666 = {1{`RANDOM}};
  _T_1010_im = _RAND_1666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1667 = {1{`RANDOM}};
  _T_1011_re = _RAND_1667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1668 = {1{`RANDOM}};
  _T_1011_im = _RAND_1668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1669 = {1{`RANDOM}};
  _T_1012_re = _RAND_1669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1670 = {1{`RANDOM}};
  _T_1012_im = _RAND_1670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1671 = {1{`RANDOM}};
  _T_1013_re = _RAND_1671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1672 = {1{`RANDOM}};
  _T_1013_im = _RAND_1672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1673 = {1{`RANDOM}};
  _T_1014_re = _RAND_1673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1674 = {1{`RANDOM}};
  _T_1014_im = _RAND_1674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1675 = {1{`RANDOM}};
  _T_1015_re = _RAND_1675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1676 = {1{`RANDOM}};
  _T_1015_im = _RAND_1676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1677 = {1{`RANDOM}};
  _T_1016_re = _RAND_1677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1678 = {1{`RANDOM}};
  _T_1016_im = _RAND_1678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1679 = {1{`RANDOM}};
  _T_1017_re = _RAND_1679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1680 = {1{`RANDOM}};
  _T_1017_im = _RAND_1680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1681 = {1{`RANDOM}};
  _T_1018_re = _RAND_1681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1682 = {1{`RANDOM}};
  _T_1018_im = _RAND_1682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1683 = {1{`RANDOM}};
  _T_1019_re = _RAND_1683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1684 = {1{`RANDOM}};
  _T_1019_im = _RAND_1684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1685 = {1{`RANDOM}};
  _T_1020_re = _RAND_1685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1686 = {1{`RANDOM}};
  _T_1020_im = _RAND_1686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1687 = {1{`RANDOM}};
  _T_1021_re = _RAND_1687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1688 = {1{`RANDOM}};
  _T_1021_im = _RAND_1688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1689 = {1{`RANDOM}};
  _T_1022_re = _RAND_1689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1690 = {1{`RANDOM}};
  _T_1022_im = _RAND_1690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1691 = {1{`RANDOM}};
  _T_1023_re = _RAND_1691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1692 = {1{`RANDOM}};
  _T_1023_im = _RAND_1692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1693 = {1{`RANDOM}};
  _T_1024_re = _RAND_1693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1694 = {1{`RANDOM}};
  _T_1024_im = _RAND_1694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1695 = {1{`RANDOM}};
  _T_1025_re = _RAND_1695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1696 = {1{`RANDOM}};
  _T_1025_im = _RAND_1696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1697 = {1{`RANDOM}};
  _T_1026_re = _RAND_1697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1698 = {1{`RANDOM}};
  _T_1026_im = _RAND_1698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1699 = {1{`RANDOM}};
  _T_1027_re = _RAND_1699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1700 = {1{`RANDOM}};
  _T_1027_im = _RAND_1700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1701 = {1{`RANDOM}};
  _T_1028_re = _RAND_1701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1702 = {1{`RANDOM}};
  _T_1028_im = _RAND_1702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1703 = {1{`RANDOM}};
  _T_1029_re = _RAND_1703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1704 = {1{`RANDOM}};
  _T_1029_im = _RAND_1704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1705 = {1{`RANDOM}};
  _T_1030_re = _RAND_1705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1706 = {1{`RANDOM}};
  _T_1030_im = _RAND_1706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1707 = {1{`RANDOM}};
  _T_1031_re = _RAND_1707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1708 = {1{`RANDOM}};
  _T_1031_im = _RAND_1708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1709 = {1{`RANDOM}};
  _T_1032_re = _RAND_1709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1710 = {1{`RANDOM}};
  _T_1032_im = _RAND_1710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1711 = {1{`RANDOM}};
  _T_1033_re = _RAND_1711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1712 = {1{`RANDOM}};
  _T_1033_im = _RAND_1712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1713 = {1{`RANDOM}};
  _T_1034_re = _RAND_1713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1714 = {1{`RANDOM}};
  _T_1034_im = _RAND_1714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1715 = {1{`RANDOM}};
  _T_1035_re = _RAND_1715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1716 = {1{`RANDOM}};
  _T_1035_im = _RAND_1716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1717 = {1{`RANDOM}};
  _T_1036_re = _RAND_1717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1718 = {1{`RANDOM}};
  _T_1036_im = _RAND_1718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1719 = {1{`RANDOM}};
  _T_1037_re = _RAND_1719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1720 = {1{`RANDOM}};
  _T_1037_im = _RAND_1720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1721 = {1{`RANDOM}};
  _T_1038_re = _RAND_1721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1722 = {1{`RANDOM}};
  _T_1038_im = _RAND_1722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1723 = {1{`RANDOM}};
  _T_1039_re = _RAND_1723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1724 = {1{`RANDOM}};
  _T_1039_im = _RAND_1724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1725 = {1{`RANDOM}};
  _T_1040_re = _RAND_1725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1726 = {1{`RANDOM}};
  _T_1040_im = _RAND_1726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1727 = {1{`RANDOM}};
  _T_1041_re = _RAND_1727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1728 = {1{`RANDOM}};
  _T_1041_im = _RAND_1728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1729 = {1{`RANDOM}};
  _T_1042_re = _RAND_1729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1730 = {1{`RANDOM}};
  _T_1042_im = _RAND_1730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1731 = {1{`RANDOM}};
  _T_1043_re = _RAND_1731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1732 = {1{`RANDOM}};
  _T_1043_im = _RAND_1732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1733 = {1{`RANDOM}};
  _T_1044_re = _RAND_1733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1734 = {1{`RANDOM}};
  _T_1044_im = _RAND_1734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1735 = {1{`RANDOM}};
  _T_1045_re = _RAND_1735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1736 = {1{`RANDOM}};
  _T_1045_im = _RAND_1736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1737 = {1{`RANDOM}};
  _T_1046_re = _RAND_1737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1738 = {1{`RANDOM}};
  _T_1046_im = _RAND_1738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1739 = {1{`RANDOM}};
  _T_1047_re = _RAND_1739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1740 = {1{`RANDOM}};
  _T_1047_im = _RAND_1740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1741 = {1{`RANDOM}};
  _T_1048_re = _RAND_1741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1742 = {1{`RANDOM}};
  _T_1048_im = _RAND_1742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1743 = {1{`RANDOM}};
  _T_1049_re = _RAND_1743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1744 = {1{`RANDOM}};
  _T_1049_im = _RAND_1744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1745 = {1{`RANDOM}};
  _T_1050_re = _RAND_1745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1746 = {1{`RANDOM}};
  _T_1050_im = _RAND_1746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1747 = {1{`RANDOM}};
  _T_1051_re = _RAND_1747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1748 = {1{`RANDOM}};
  _T_1051_im = _RAND_1748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1749 = {1{`RANDOM}};
  _T_1052_re = _RAND_1749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1750 = {1{`RANDOM}};
  _T_1052_im = _RAND_1750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1751 = {1{`RANDOM}};
  _T_1053_re = _RAND_1751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1752 = {1{`RANDOM}};
  _T_1053_im = _RAND_1752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1753 = {1{`RANDOM}};
  _T_1054_re = _RAND_1753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1754 = {1{`RANDOM}};
  _T_1054_im = _RAND_1754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1755 = {1{`RANDOM}};
  _T_1055_re = _RAND_1755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1756 = {1{`RANDOM}};
  _T_1055_im = _RAND_1756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1757 = {1{`RANDOM}};
  _T_1056_re = _RAND_1757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1758 = {1{`RANDOM}};
  _T_1056_im = _RAND_1758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1759 = {1{`RANDOM}};
  _T_1057_re = _RAND_1759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1760 = {1{`RANDOM}};
  _T_1057_im = _RAND_1760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1761 = {1{`RANDOM}};
  _T_1058_re = _RAND_1761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1762 = {1{`RANDOM}};
  _T_1058_im = _RAND_1762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1763 = {1{`RANDOM}};
  _T_1059_re = _RAND_1763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1764 = {1{`RANDOM}};
  _T_1059_im = _RAND_1764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1765 = {1{`RANDOM}};
  _T_1060_re = _RAND_1765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1766 = {1{`RANDOM}};
  _T_1060_im = _RAND_1766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1767 = {1{`RANDOM}};
  _T_1061_re = _RAND_1767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1768 = {1{`RANDOM}};
  _T_1061_im = _RAND_1768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1769 = {1{`RANDOM}};
  _T_1062_re = _RAND_1769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1770 = {1{`RANDOM}};
  _T_1062_im = _RAND_1770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1771 = {1{`RANDOM}};
  _T_1063_re = _RAND_1771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1772 = {1{`RANDOM}};
  _T_1063_im = _RAND_1772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1773 = {1{`RANDOM}};
  _T_1064_re = _RAND_1773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1774 = {1{`RANDOM}};
  _T_1064_im = _RAND_1774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1775 = {1{`RANDOM}};
  _T_1065_re = _RAND_1775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1776 = {1{`RANDOM}};
  _T_1065_im = _RAND_1776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1777 = {1{`RANDOM}};
  _T_1066_re = _RAND_1777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1778 = {1{`RANDOM}};
  _T_1066_im = _RAND_1778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1779 = {1{`RANDOM}};
  _T_1067_re = _RAND_1779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1780 = {1{`RANDOM}};
  _T_1067_im = _RAND_1780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1781 = {1{`RANDOM}};
  _T_1068_re = _RAND_1781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1782 = {1{`RANDOM}};
  _T_1068_im = _RAND_1782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1783 = {1{`RANDOM}};
  _T_1069_re = _RAND_1783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1784 = {1{`RANDOM}};
  _T_1069_im = _RAND_1784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1785 = {1{`RANDOM}};
  _T_1070_re = _RAND_1785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1786 = {1{`RANDOM}};
  _T_1070_im = _RAND_1786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1787 = {1{`RANDOM}};
  _T_1071_re = _RAND_1787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1788 = {1{`RANDOM}};
  _T_1071_im = _RAND_1788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1789 = {1{`RANDOM}};
  _T_1072_re = _RAND_1789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1790 = {1{`RANDOM}};
  _T_1072_im = _RAND_1790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1791 = {1{`RANDOM}};
  _T_1073_re = _RAND_1791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1792 = {1{`RANDOM}};
  _T_1073_im = _RAND_1792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1793 = {1{`RANDOM}};
  _T_1074_re = _RAND_1793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1794 = {1{`RANDOM}};
  _T_1074_im = _RAND_1794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1795 = {1{`RANDOM}};
  _T_1075_re = _RAND_1795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1796 = {1{`RANDOM}};
  _T_1075_im = _RAND_1796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1797 = {1{`RANDOM}};
  _T_1076_re = _RAND_1797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1798 = {1{`RANDOM}};
  _T_1076_im = _RAND_1798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1799 = {1{`RANDOM}};
  _T_1077_re = _RAND_1799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1800 = {1{`RANDOM}};
  _T_1077_im = _RAND_1800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1801 = {1{`RANDOM}};
  _T_1078_re = _RAND_1801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1802 = {1{`RANDOM}};
  _T_1078_im = _RAND_1802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1803 = {1{`RANDOM}};
  _T_1079_re = _RAND_1803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1804 = {1{`RANDOM}};
  _T_1079_im = _RAND_1804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1805 = {1{`RANDOM}};
  _T_1080_re = _RAND_1805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1806 = {1{`RANDOM}};
  _T_1080_im = _RAND_1806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1807 = {1{`RANDOM}};
  _T_1081_re = _RAND_1807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1808 = {1{`RANDOM}};
  _T_1081_im = _RAND_1808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1809 = {1{`RANDOM}};
  _T_1082_re = _RAND_1809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1810 = {1{`RANDOM}};
  _T_1082_im = _RAND_1810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1811 = {1{`RANDOM}};
  _T_1083_re = _RAND_1811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1812 = {1{`RANDOM}};
  _T_1083_im = _RAND_1812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1813 = {1{`RANDOM}};
  _T_1084_re = _RAND_1813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1814 = {1{`RANDOM}};
  _T_1084_im = _RAND_1814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1815 = {1{`RANDOM}};
  _T_1085_re = _RAND_1815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1816 = {1{`RANDOM}};
  _T_1085_im = _RAND_1816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1817 = {1{`RANDOM}};
  _T_1086_re = _RAND_1817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1818 = {1{`RANDOM}};
  _T_1086_im = _RAND_1818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1819 = {1{`RANDOM}};
  _T_1087_re = _RAND_1819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1820 = {1{`RANDOM}};
  _T_1087_im = _RAND_1820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1821 = {1{`RANDOM}};
  _T_1088_re = _RAND_1821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1822 = {1{`RANDOM}};
  _T_1088_im = _RAND_1822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1823 = {1{`RANDOM}};
  _T_1089_re = _RAND_1823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1824 = {1{`RANDOM}};
  _T_1089_im = _RAND_1824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1825 = {1{`RANDOM}};
  _T_1090_re = _RAND_1825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1826 = {1{`RANDOM}};
  _T_1090_im = _RAND_1826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1827 = {1{`RANDOM}};
  _T_1091_re = _RAND_1827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1828 = {1{`RANDOM}};
  _T_1091_im = _RAND_1828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1829 = {1{`RANDOM}};
  _T_1092_re = _RAND_1829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1830 = {1{`RANDOM}};
  _T_1092_im = _RAND_1830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1831 = {1{`RANDOM}};
  _T_1093_re = _RAND_1831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1832 = {1{`RANDOM}};
  _T_1093_im = _RAND_1832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1833 = {1{`RANDOM}};
  _T_1094_re = _RAND_1833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1834 = {1{`RANDOM}};
  _T_1094_im = _RAND_1834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1835 = {1{`RANDOM}};
  _T_1095_re = _RAND_1835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1836 = {1{`RANDOM}};
  _T_1095_im = _RAND_1836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1837 = {1{`RANDOM}};
  _T_1096_re = _RAND_1837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1838 = {1{`RANDOM}};
  _T_1096_im = _RAND_1838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1839 = {1{`RANDOM}};
  _T_1097_re = _RAND_1839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1840 = {1{`RANDOM}};
  _T_1097_im = _RAND_1840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1841 = {1{`RANDOM}};
  _T_1098_re = _RAND_1841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1842 = {1{`RANDOM}};
  _T_1098_im = _RAND_1842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1843 = {1{`RANDOM}};
  _T_1099_re = _RAND_1843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1844 = {1{`RANDOM}};
  _T_1099_im = _RAND_1844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1845 = {1{`RANDOM}};
  _T_1100_re = _RAND_1845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1846 = {1{`RANDOM}};
  _T_1100_im = _RAND_1846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1847 = {1{`RANDOM}};
  _T_1101_re = _RAND_1847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1848 = {1{`RANDOM}};
  _T_1101_im = _RAND_1848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1849 = {1{`RANDOM}};
  _T_1102_re = _RAND_1849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1850 = {1{`RANDOM}};
  _T_1102_im = _RAND_1850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1851 = {1{`RANDOM}};
  _T_1103_re = _RAND_1851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1852 = {1{`RANDOM}};
  _T_1103_im = _RAND_1852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1853 = {1{`RANDOM}};
  _T_1104_re = _RAND_1853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1854 = {1{`RANDOM}};
  _T_1104_im = _RAND_1854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1855 = {1{`RANDOM}};
  _T_1105_re = _RAND_1855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1856 = {1{`RANDOM}};
  _T_1105_im = _RAND_1856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1857 = {1{`RANDOM}};
  _T_1106_re = _RAND_1857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1858 = {1{`RANDOM}};
  _T_1106_im = _RAND_1858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1859 = {1{`RANDOM}};
  _T_1107_re = _RAND_1859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1860 = {1{`RANDOM}};
  _T_1107_im = _RAND_1860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1861 = {1{`RANDOM}};
  _T_1108_re = _RAND_1861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1862 = {1{`RANDOM}};
  _T_1108_im = _RAND_1862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1863 = {1{`RANDOM}};
  _T_1109_re = _RAND_1863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1864 = {1{`RANDOM}};
  _T_1109_im = _RAND_1864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1865 = {1{`RANDOM}};
  _T_1110_re = _RAND_1865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1866 = {1{`RANDOM}};
  _T_1110_im = _RAND_1866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1867 = {1{`RANDOM}};
  _T_1111_re = _RAND_1867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1868 = {1{`RANDOM}};
  _T_1111_im = _RAND_1868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1869 = {1{`RANDOM}};
  _T_1112_re = _RAND_1869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1870 = {1{`RANDOM}};
  _T_1112_im = _RAND_1870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1871 = {1{`RANDOM}};
  _T_1113_re = _RAND_1871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1872 = {1{`RANDOM}};
  _T_1113_im = _RAND_1872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1873 = {1{`RANDOM}};
  _T_1114_re = _RAND_1873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1874 = {1{`RANDOM}};
  _T_1114_im = _RAND_1874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1875 = {1{`RANDOM}};
  _T_1115_re = _RAND_1875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1876 = {1{`RANDOM}};
  _T_1115_im = _RAND_1876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1877 = {1{`RANDOM}};
  _T_1116_re = _RAND_1877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1878 = {1{`RANDOM}};
  _T_1116_im = _RAND_1878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1879 = {1{`RANDOM}};
  _T_1117_re = _RAND_1879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1880 = {1{`RANDOM}};
  _T_1117_im = _RAND_1880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1881 = {1{`RANDOM}};
  _T_1118_re = _RAND_1881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1882 = {1{`RANDOM}};
  _T_1118_im = _RAND_1882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1883 = {1{`RANDOM}};
  _T_1119_re = _RAND_1883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1884 = {1{`RANDOM}};
  _T_1119_im = _RAND_1884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1885 = {1{`RANDOM}};
  _T_1120_re = _RAND_1885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1886 = {1{`RANDOM}};
  _T_1120_im = _RAND_1886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1887 = {1{`RANDOM}};
  _T_1121_re = _RAND_1887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1888 = {1{`RANDOM}};
  _T_1121_im = _RAND_1888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1889 = {1{`RANDOM}};
  _T_1122_re = _RAND_1889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1890 = {1{`RANDOM}};
  _T_1122_im = _RAND_1890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1891 = {1{`RANDOM}};
  _T_1123_re = _RAND_1891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1892 = {1{`RANDOM}};
  _T_1123_im = _RAND_1892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1893 = {1{`RANDOM}};
  _T_1124_re = _RAND_1893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1894 = {1{`RANDOM}};
  _T_1124_im = _RAND_1894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1895 = {1{`RANDOM}};
  _T_1125_re = _RAND_1895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1896 = {1{`RANDOM}};
  _T_1125_im = _RAND_1896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1897 = {1{`RANDOM}};
  _T_1126_re = _RAND_1897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1898 = {1{`RANDOM}};
  _T_1126_im = _RAND_1898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1899 = {1{`RANDOM}};
  _T_1127_re = _RAND_1899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1900 = {1{`RANDOM}};
  _T_1127_im = _RAND_1900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1901 = {1{`RANDOM}};
  _T_1128_re = _RAND_1901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1902 = {1{`RANDOM}};
  _T_1128_im = _RAND_1902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1903 = {1{`RANDOM}};
  _T_1129_re = _RAND_1903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1904 = {1{`RANDOM}};
  _T_1129_im = _RAND_1904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1905 = {1{`RANDOM}};
  _T_1130_re = _RAND_1905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1906 = {1{`RANDOM}};
  _T_1130_im = _RAND_1906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1907 = {1{`RANDOM}};
  _T_1131_re = _RAND_1907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1908 = {1{`RANDOM}};
  _T_1131_im = _RAND_1908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1909 = {1{`RANDOM}};
  _T_1132_re = _RAND_1909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1910 = {1{`RANDOM}};
  _T_1132_im = _RAND_1910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1911 = {1{`RANDOM}};
  _T_1133_re = _RAND_1911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1912 = {1{`RANDOM}};
  _T_1133_im = _RAND_1912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1913 = {1{`RANDOM}};
  _T_1134_re = _RAND_1913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1914 = {1{`RANDOM}};
  _T_1134_im = _RAND_1914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1915 = {1{`RANDOM}};
  _T_1135_re = _RAND_1915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1916 = {1{`RANDOM}};
  _T_1135_im = _RAND_1916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1917 = {1{`RANDOM}};
  _T_1136_re = _RAND_1917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1918 = {1{`RANDOM}};
  _T_1136_im = _RAND_1918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1919 = {1{`RANDOM}};
  _T_1137_re = _RAND_1919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1920 = {1{`RANDOM}};
  _T_1137_im = _RAND_1920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1921 = {1{`RANDOM}};
  _T_1138_re = _RAND_1921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1922 = {1{`RANDOM}};
  _T_1138_im = _RAND_1922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1923 = {1{`RANDOM}};
  _T_1139_re = _RAND_1923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1924 = {1{`RANDOM}};
  _T_1139_im = _RAND_1924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1925 = {1{`RANDOM}};
  _T_1140_re = _RAND_1925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1926 = {1{`RANDOM}};
  _T_1140_im = _RAND_1926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1927 = {1{`RANDOM}};
  _T_1141_re = _RAND_1927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1928 = {1{`RANDOM}};
  _T_1141_im = _RAND_1928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1929 = {1{`RANDOM}};
  _T_1142_re = _RAND_1929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1930 = {1{`RANDOM}};
  _T_1142_im = _RAND_1930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1931 = {1{`RANDOM}};
  _T_1143_re = _RAND_1931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1932 = {1{`RANDOM}};
  _T_1143_im = _RAND_1932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1933 = {1{`RANDOM}};
  _T_1144_re = _RAND_1933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1934 = {1{`RANDOM}};
  _T_1144_im = _RAND_1934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1935 = {1{`RANDOM}};
  _T_1145_re = _RAND_1935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1936 = {1{`RANDOM}};
  _T_1145_im = _RAND_1936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1937 = {1{`RANDOM}};
  _T_1146_re = _RAND_1937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1938 = {1{`RANDOM}};
  _T_1146_im = _RAND_1938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1939 = {1{`RANDOM}};
  _T_1147_re = _RAND_1939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1940 = {1{`RANDOM}};
  _T_1147_im = _RAND_1940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1941 = {1{`RANDOM}};
  _T_1148_re = _RAND_1941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1942 = {1{`RANDOM}};
  _T_1148_im = _RAND_1942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1943 = {1{`RANDOM}};
  _T_1149_re = _RAND_1943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1944 = {1{`RANDOM}};
  _T_1149_im = _RAND_1944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1945 = {1{`RANDOM}};
  _T_1150_re = _RAND_1945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1946 = {1{`RANDOM}};
  _T_1150_im = _RAND_1946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1947 = {1{`RANDOM}};
  _T_1151_re = _RAND_1947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1948 = {1{`RANDOM}};
  _T_1151_im = _RAND_1948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1949 = {1{`RANDOM}};
  _T_1152_re = _RAND_1949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1950 = {1{`RANDOM}};
  _T_1152_im = _RAND_1950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1951 = {1{`RANDOM}};
  _T_1153_re = _RAND_1951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1952 = {1{`RANDOM}};
  _T_1153_im = _RAND_1952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1953 = {1{`RANDOM}};
  _T_1154_re = _RAND_1953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1954 = {1{`RANDOM}};
  _T_1154_im = _RAND_1954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1955 = {1{`RANDOM}};
  _T_1155_re = _RAND_1955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1956 = {1{`RANDOM}};
  _T_1155_im = _RAND_1956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1957 = {1{`RANDOM}};
  _T_1156_re = _RAND_1957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1958 = {1{`RANDOM}};
  _T_1156_im = _RAND_1958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1959 = {1{`RANDOM}};
  _T_1157_re = _RAND_1959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1960 = {1{`RANDOM}};
  _T_1157_im = _RAND_1960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1961 = {1{`RANDOM}};
  _T_1158_re = _RAND_1961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1962 = {1{`RANDOM}};
  _T_1158_im = _RAND_1962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1963 = {1{`RANDOM}};
  _T_1159_re = _RAND_1963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1964 = {1{`RANDOM}};
  _T_1159_im = _RAND_1964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1965 = {1{`RANDOM}};
  _T_1160_re = _RAND_1965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1966 = {1{`RANDOM}};
  _T_1160_im = _RAND_1966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1967 = {1{`RANDOM}};
  _T_1161_re = _RAND_1967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1968 = {1{`RANDOM}};
  _T_1161_im = _RAND_1968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1969 = {1{`RANDOM}};
  _T_1162_re = _RAND_1969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1970 = {1{`RANDOM}};
  _T_1162_im = _RAND_1970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1971 = {1{`RANDOM}};
  _T_1163_re = _RAND_1971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1972 = {1{`RANDOM}};
  _T_1163_im = _RAND_1972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1973 = {1{`RANDOM}};
  _T_1164_re = _RAND_1973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1974 = {1{`RANDOM}};
  _T_1164_im = _RAND_1974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1975 = {1{`RANDOM}};
  _T_1165_re = _RAND_1975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1976 = {1{`RANDOM}};
  _T_1165_im = _RAND_1976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1977 = {1{`RANDOM}};
  _T_1166_re = _RAND_1977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1978 = {1{`RANDOM}};
  _T_1166_im = _RAND_1978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1979 = {1{`RANDOM}};
  _T_1167_re = _RAND_1979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1980 = {1{`RANDOM}};
  _T_1167_im = _RAND_1980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1981 = {1{`RANDOM}};
  _T_1168_re = _RAND_1981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1982 = {1{`RANDOM}};
  _T_1168_im = _RAND_1982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1983 = {1{`RANDOM}};
  _T_1169_re = _RAND_1983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1984 = {1{`RANDOM}};
  _T_1169_im = _RAND_1984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1985 = {1{`RANDOM}};
  _T_1170_re = _RAND_1985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1986 = {1{`RANDOM}};
  _T_1170_im = _RAND_1986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1987 = {1{`RANDOM}};
  _T_1171_re = _RAND_1987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1988 = {1{`RANDOM}};
  _T_1171_im = _RAND_1988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1989 = {1{`RANDOM}};
  _T_1172_re = _RAND_1989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1990 = {1{`RANDOM}};
  _T_1172_im = _RAND_1990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1991 = {1{`RANDOM}};
  _T_1173_re = _RAND_1991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1992 = {1{`RANDOM}};
  _T_1173_im = _RAND_1992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1993 = {1{`RANDOM}};
  _T_1174_re = _RAND_1993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1994 = {1{`RANDOM}};
  _T_1174_im = _RAND_1994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1995 = {1{`RANDOM}};
  _T_1175_re = _RAND_1995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1996 = {1{`RANDOM}};
  _T_1175_im = _RAND_1996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1997 = {1{`RANDOM}};
  _T_1176_re = _RAND_1997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1998 = {1{`RANDOM}};
  _T_1176_im = _RAND_1998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1999 = {1{`RANDOM}};
  _T_1177_re = _RAND_1999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2000 = {1{`RANDOM}};
  _T_1177_im = _RAND_2000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2001 = {1{`RANDOM}};
  _T_1178_re = _RAND_2001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2002 = {1{`RANDOM}};
  _T_1178_im = _RAND_2002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2003 = {1{`RANDOM}};
  _T_1179_re = _RAND_2003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2004 = {1{`RANDOM}};
  _T_1179_im = _RAND_2004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2005 = {1{`RANDOM}};
  _T_1180_re = _RAND_2005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2006 = {1{`RANDOM}};
  _T_1180_im = _RAND_2006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2007 = {1{`RANDOM}};
  _T_1181_re = _RAND_2007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2008 = {1{`RANDOM}};
  _T_1181_im = _RAND_2008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2009 = {1{`RANDOM}};
  _T_1182_re = _RAND_2009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2010 = {1{`RANDOM}};
  _T_1182_im = _RAND_2010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2011 = {1{`RANDOM}};
  _T_1183_re = _RAND_2011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2012 = {1{`RANDOM}};
  _T_1183_im = _RAND_2012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2013 = {1{`RANDOM}};
  _T_1184_re = _RAND_2013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2014 = {1{`RANDOM}};
  _T_1184_im = _RAND_2014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2015 = {1{`RANDOM}};
  _T_1185_re = _RAND_2015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2016 = {1{`RANDOM}};
  _T_1185_im = _RAND_2016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2017 = {1{`RANDOM}};
  _T_1186_re = _RAND_2017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2018 = {1{`RANDOM}};
  _T_1186_im = _RAND_2018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2019 = {1{`RANDOM}};
  _T_1187_re = _RAND_2019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2020 = {1{`RANDOM}};
  _T_1187_im = _RAND_2020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2021 = {1{`RANDOM}};
  _T_1188_re = _RAND_2021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2022 = {1{`RANDOM}};
  _T_1188_im = _RAND_2022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2023 = {1{`RANDOM}};
  _T_1189_re = _RAND_2023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2024 = {1{`RANDOM}};
  _T_1189_im = _RAND_2024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2025 = {1{`RANDOM}};
  _T_1190_re = _RAND_2025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2026 = {1{`RANDOM}};
  _T_1190_im = _RAND_2026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2027 = {1{`RANDOM}};
  _T_1191_re = _RAND_2027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2028 = {1{`RANDOM}};
  _T_1191_im = _RAND_2028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2029 = {1{`RANDOM}};
  _T_1192_re = _RAND_2029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2030 = {1{`RANDOM}};
  _T_1192_im = _RAND_2030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2031 = {1{`RANDOM}};
  _T_1193_re = _RAND_2031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2032 = {1{`RANDOM}};
  _T_1193_im = _RAND_2032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2033 = {1{`RANDOM}};
  _T_1194_re = _RAND_2033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2034 = {1{`RANDOM}};
  _T_1194_im = _RAND_2034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2035 = {1{`RANDOM}};
  _T_1195_re = _RAND_2035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2036 = {1{`RANDOM}};
  _T_1195_im = _RAND_2036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2037 = {1{`RANDOM}};
  _T_1196_re = _RAND_2037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2038 = {1{`RANDOM}};
  _T_1196_im = _RAND_2038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2039 = {1{`RANDOM}};
  _T_1197_re = _RAND_2039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2040 = {1{`RANDOM}};
  _T_1197_im = _RAND_2040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2041 = {1{`RANDOM}};
  _T_1198_re = _RAND_2041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2042 = {1{`RANDOM}};
  _T_1198_im = _RAND_2042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2043 = {1{`RANDOM}};
  _T_1199_re = _RAND_2043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2044 = {1{`RANDOM}};
  _T_1199_im = _RAND_2044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2045 = {1{`RANDOM}};
  _T_1200_re = _RAND_2045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2046 = {1{`RANDOM}};
  _T_1200_im = _RAND_2046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2047 = {1{`RANDOM}};
  _T_1201_re = _RAND_2047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2048 = {1{`RANDOM}};
  _T_1201_im = _RAND_2048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2049 = {1{`RANDOM}};
  _T_1202_re = _RAND_2049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2050 = {1{`RANDOM}};
  _T_1202_im = _RAND_2050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2051 = {1{`RANDOM}};
  _T_1203_re = _RAND_2051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2052 = {1{`RANDOM}};
  _T_1203_im = _RAND_2052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2053 = {1{`RANDOM}};
  _T_1204_re = _RAND_2053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2054 = {1{`RANDOM}};
  _T_1204_im = _RAND_2054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2055 = {1{`RANDOM}};
  _T_1207_re = _RAND_2055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2056 = {1{`RANDOM}};
  _T_1207_im = _RAND_2056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2057 = {1{`RANDOM}};
  _T_1208_re = _RAND_2057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2058 = {1{`RANDOM}};
  _T_1208_im = _RAND_2058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2059 = {1{`RANDOM}};
  _T_1209_re = _RAND_2059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2060 = {1{`RANDOM}};
  _T_1209_im = _RAND_2060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2061 = {1{`RANDOM}};
  _T_1210_re = _RAND_2061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2062 = {1{`RANDOM}};
  _T_1210_im = _RAND_2062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2063 = {1{`RANDOM}};
  _T_1211_re = _RAND_2063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2064 = {1{`RANDOM}};
  _T_1211_im = _RAND_2064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2065 = {1{`RANDOM}};
  _T_1212_re = _RAND_2065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2066 = {1{`RANDOM}};
  _T_1212_im = _RAND_2066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2067 = {1{`RANDOM}};
  _T_1213_re = _RAND_2067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2068 = {1{`RANDOM}};
  _T_1213_im = _RAND_2068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2069 = {1{`RANDOM}};
  _T_1214_re = _RAND_2069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2070 = {1{`RANDOM}};
  _T_1214_im = _RAND_2070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2071 = {1{`RANDOM}};
  _T_1215_re = _RAND_2071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2072 = {1{`RANDOM}};
  _T_1215_im = _RAND_2072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2073 = {1{`RANDOM}};
  _T_1216_re = _RAND_2073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2074 = {1{`RANDOM}};
  _T_1216_im = _RAND_2074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2075 = {1{`RANDOM}};
  _T_1217_re = _RAND_2075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2076 = {1{`RANDOM}};
  _T_1217_im = _RAND_2076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2077 = {1{`RANDOM}};
  _T_1218_re = _RAND_2077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2078 = {1{`RANDOM}};
  _T_1218_im = _RAND_2078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2079 = {1{`RANDOM}};
  _T_1219_re = _RAND_2079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2080 = {1{`RANDOM}};
  _T_1219_im = _RAND_2080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2081 = {1{`RANDOM}};
  _T_1220_re = _RAND_2081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2082 = {1{`RANDOM}};
  _T_1220_im = _RAND_2082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2083 = {1{`RANDOM}};
  _T_1221_re = _RAND_2083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2084 = {1{`RANDOM}};
  _T_1221_im = _RAND_2084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2085 = {1{`RANDOM}};
  _T_1222_re = _RAND_2085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2086 = {1{`RANDOM}};
  _T_1222_im = _RAND_2086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2087 = {1{`RANDOM}};
  _T_1223_re = _RAND_2087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2088 = {1{`RANDOM}};
  _T_1223_im = _RAND_2088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2089 = {1{`RANDOM}};
  _T_1224_re = _RAND_2089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2090 = {1{`RANDOM}};
  _T_1224_im = _RAND_2090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2091 = {1{`RANDOM}};
  _T_1225_re = _RAND_2091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2092 = {1{`RANDOM}};
  _T_1225_im = _RAND_2092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2093 = {1{`RANDOM}};
  _T_1226_re = _RAND_2093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2094 = {1{`RANDOM}};
  _T_1226_im = _RAND_2094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2095 = {1{`RANDOM}};
  _T_1227_re = _RAND_2095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2096 = {1{`RANDOM}};
  _T_1227_im = _RAND_2096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2097 = {1{`RANDOM}};
  _T_1228_re = _RAND_2097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2098 = {1{`RANDOM}};
  _T_1228_im = _RAND_2098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2099 = {1{`RANDOM}};
  _T_1229_re = _RAND_2099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2100 = {1{`RANDOM}};
  _T_1229_im = _RAND_2100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2101 = {1{`RANDOM}};
  _T_1230_re = _RAND_2101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2102 = {1{`RANDOM}};
  _T_1230_im = _RAND_2102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2103 = {1{`RANDOM}};
  _T_1231_re = _RAND_2103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2104 = {1{`RANDOM}};
  _T_1231_im = _RAND_2104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2105 = {1{`RANDOM}};
  _T_1232_re = _RAND_2105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2106 = {1{`RANDOM}};
  _T_1232_im = _RAND_2106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2107 = {1{`RANDOM}};
  _T_1233_re = _RAND_2107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2108 = {1{`RANDOM}};
  _T_1233_im = _RAND_2108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2109 = {1{`RANDOM}};
  _T_1234_re = _RAND_2109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2110 = {1{`RANDOM}};
  _T_1234_im = _RAND_2110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2111 = {1{`RANDOM}};
  _T_1235_re = _RAND_2111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2112 = {1{`RANDOM}};
  _T_1235_im = _RAND_2112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2113 = {1{`RANDOM}};
  _T_1236_re = _RAND_2113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2114 = {1{`RANDOM}};
  _T_1236_im = _RAND_2114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2115 = {1{`RANDOM}};
  _T_1237_re = _RAND_2115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2116 = {1{`RANDOM}};
  _T_1237_im = _RAND_2116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2117 = {1{`RANDOM}};
  _T_1238_re = _RAND_2117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2118 = {1{`RANDOM}};
  _T_1238_im = _RAND_2118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2119 = {1{`RANDOM}};
  _T_1239_re = _RAND_2119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2120 = {1{`RANDOM}};
  _T_1239_im = _RAND_2120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2121 = {1{`RANDOM}};
  _T_1240_re = _RAND_2121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2122 = {1{`RANDOM}};
  _T_1240_im = _RAND_2122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2123 = {1{`RANDOM}};
  _T_1241_re = _RAND_2123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2124 = {1{`RANDOM}};
  _T_1241_im = _RAND_2124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2125 = {1{`RANDOM}};
  _T_1242_re = _RAND_2125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2126 = {1{`RANDOM}};
  _T_1242_im = _RAND_2126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2127 = {1{`RANDOM}};
  _T_1243_re = _RAND_2127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2128 = {1{`RANDOM}};
  _T_1243_im = _RAND_2128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2129 = {1{`RANDOM}};
  _T_1244_re = _RAND_2129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2130 = {1{`RANDOM}};
  _T_1244_im = _RAND_2130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2131 = {1{`RANDOM}};
  _T_1245_re = _RAND_2131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2132 = {1{`RANDOM}};
  _T_1245_im = _RAND_2132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2133 = {1{`RANDOM}};
  _T_1246_re = _RAND_2133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2134 = {1{`RANDOM}};
  _T_1246_im = _RAND_2134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2135 = {1{`RANDOM}};
  _T_1247_re = _RAND_2135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2136 = {1{`RANDOM}};
  _T_1247_im = _RAND_2136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2137 = {1{`RANDOM}};
  _T_1248_re = _RAND_2137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2138 = {1{`RANDOM}};
  _T_1248_im = _RAND_2138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2139 = {1{`RANDOM}};
  _T_1249_re = _RAND_2139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2140 = {1{`RANDOM}};
  _T_1249_im = _RAND_2140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2141 = {1{`RANDOM}};
  _T_1250_re = _RAND_2141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2142 = {1{`RANDOM}};
  _T_1250_im = _RAND_2142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2143 = {1{`RANDOM}};
  _T_1251_re = _RAND_2143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2144 = {1{`RANDOM}};
  _T_1251_im = _RAND_2144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2145 = {1{`RANDOM}};
  _T_1252_re = _RAND_2145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2146 = {1{`RANDOM}};
  _T_1252_im = _RAND_2146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2147 = {1{`RANDOM}};
  _T_1253_re = _RAND_2147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2148 = {1{`RANDOM}};
  _T_1253_im = _RAND_2148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2149 = {1{`RANDOM}};
  _T_1254_re = _RAND_2149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2150 = {1{`RANDOM}};
  _T_1254_im = _RAND_2150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2151 = {1{`RANDOM}};
  _T_1255_re = _RAND_2151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2152 = {1{`RANDOM}};
  _T_1255_im = _RAND_2152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2153 = {1{`RANDOM}};
  _T_1256_re = _RAND_2153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2154 = {1{`RANDOM}};
  _T_1256_im = _RAND_2154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2155 = {1{`RANDOM}};
  _T_1257_re = _RAND_2155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2156 = {1{`RANDOM}};
  _T_1257_im = _RAND_2156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2157 = {1{`RANDOM}};
  _T_1258_re = _RAND_2157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2158 = {1{`RANDOM}};
  _T_1258_im = _RAND_2158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2159 = {1{`RANDOM}};
  _T_1259_re = _RAND_2159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2160 = {1{`RANDOM}};
  _T_1259_im = _RAND_2160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2161 = {1{`RANDOM}};
  _T_1260_re = _RAND_2161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2162 = {1{`RANDOM}};
  _T_1260_im = _RAND_2162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2163 = {1{`RANDOM}};
  _T_1261_re = _RAND_2163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2164 = {1{`RANDOM}};
  _T_1261_im = _RAND_2164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2165 = {1{`RANDOM}};
  _T_1262_re = _RAND_2165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2166 = {1{`RANDOM}};
  _T_1262_im = _RAND_2166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2167 = {1{`RANDOM}};
  _T_1263_re = _RAND_2167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2168 = {1{`RANDOM}};
  _T_1263_im = _RAND_2168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2169 = {1{`RANDOM}};
  _T_1264_re = _RAND_2169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2170 = {1{`RANDOM}};
  _T_1264_im = _RAND_2170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2171 = {1{`RANDOM}};
  _T_1265_re = _RAND_2171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2172 = {1{`RANDOM}};
  _T_1265_im = _RAND_2172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2173 = {1{`RANDOM}};
  _T_1266_re = _RAND_2173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2174 = {1{`RANDOM}};
  _T_1266_im = _RAND_2174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2175 = {1{`RANDOM}};
  _T_1267_re = _RAND_2175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2176 = {1{`RANDOM}};
  _T_1267_im = _RAND_2176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2177 = {1{`RANDOM}};
  _T_1268_re = _RAND_2177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2178 = {1{`RANDOM}};
  _T_1268_im = _RAND_2178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2179 = {1{`RANDOM}};
  _T_1269_re = _RAND_2179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2180 = {1{`RANDOM}};
  _T_1269_im = _RAND_2180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2181 = {1{`RANDOM}};
  _T_1270_re = _RAND_2181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2182 = {1{`RANDOM}};
  _T_1270_im = _RAND_2182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2183 = {1{`RANDOM}};
  _T_1271_re = _RAND_2183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2184 = {1{`RANDOM}};
  _T_1271_im = _RAND_2184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2185 = {1{`RANDOM}};
  _T_1272_re = _RAND_2185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2186 = {1{`RANDOM}};
  _T_1272_im = _RAND_2186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2187 = {1{`RANDOM}};
  _T_1273_re = _RAND_2187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2188 = {1{`RANDOM}};
  _T_1273_im = _RAND_2188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2189 = {1{`RANDOM}};
  _T_1274_re = _RAND_2189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2190 = {1{`RANDOM}};
  _T_1274_im = _RAND_2190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2191 = {1{`RANDOM}};
  _T_1275_re = _RAND_2191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2192 = {1{`RANDOM}};
  _T_1275_im = _RAND_2192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2193 = {1{`RANDOM}};
  _T_1276_re = _RAND_2193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2194 = {1{`RANDOM}};
  _T_1276_im = _RAND_2194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2195 = {1{`RANDOM}};
  _T_1277_re = _RAND_2195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2196 = {1{`RANDOM}};
  _T_1277_im = _RAND_2196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2197 = {1{`RANDOM}};
  _T_1278_re = _RAND_2197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2198 = {1{`RANDOM}};
  _T_1278_im = _RAND_2198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2199 = {1{`RANDOM}};
  _T_1279_re = _RAND_2199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2200 = {1{`RANDOM}};
  _T_1279_im = _RAND_2200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2201 = {1{`RANDOM}};
  _T_1280_re = _RAND_2201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2202 = {1{`RANDOM}};
  _T_1280_im = _RAND_2202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2203 = {1{`RANDOM}};
  _T_1281_re = _RAND_2203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2204 = {1{`RANDOM}};
  _T_1281_im = _RAND_2204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2205 = {1{`RANDOM}};
  _T_1282_re = _RAND_2205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2206 = {1{`RANDOM}};
  _T_1282_im = _RAND_2206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2207 = {1{`RANDOM}};
  _T_1283_re = _RAND_2207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2208 = {1{`RANDOM}};
  _T_1283_im = _RAND_2208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2209 = {1{`RANDOM}};
  _T_1284_re = _RAND_2209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2210 = {1{`RANDOM}};
  _T_1284_im = _RAND_2210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2211 = {1{`RANDOM}};
  _T_1285_re = _RAND_2211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2212 = {1{`RANDOM}};
  _T_1285_im = _RAND_2212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2213 = {1{`RANDOM}};
  _T_1286_re = _RAND_2213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2214 = {1{`RANDOM}};
  _T_1286_im = _RAND_2214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2215 = {1{`RANDOM}};
  _T_1287_re = _RAND_2215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2216 = {1{`RANDOM}};
  _T_1287_im = _RAND_2216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2217 = {1{`RANDOM}};
  _T_1288_re = _RAND_2217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2218 = {1{`RANDOM}};
  _T_1288_im = _RAND_2218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2219 = {1{`RANDOM}};
  _T_1289_re = _RAND_2219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2220 = {1{`RANDOM}};
  _T_1289_im = _RAND_2220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2221 = {1{`RANDOM}};
  _T_1290_re = _RAND_2221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2222 = {1{`RANDOM}};
  _T_1290_im = _RAND_2222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2223 = {1{`RANDOM}};
  _T_1291_re = _RAND_2223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2224 = {1{`RANDOM}};
  _T_1291_im = _RAND_2224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2225 = {1{`RANDOM}};
  _T_1292_re = _RAND_2225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2226 = {1{`RANDOM}};
  _T_1292_im = _RAND_2226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2227 = {1{`RANDOM}};
  _T_1293_re = _RAND_2227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2228 = {1{`RANDOM}};
  _T_1293_im = _RAND_2228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2229 = {1{`RANDOM}};
  _T_1294_re = _RAND_2229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2230 = {1{`RANDOM}};
  _T_1294_im = _RAND_2230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2231 = {1{`RANDOM}};
  _T_1295_re = _RAND_2231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2232 = {1{`RANDOM}};
  _T_1295_im = _RAND_2232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2233 = {1{`RANDOM}};
  _T_1296_re = _RAND_2233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2234 = {1{`RANDOM}};
  _T_1296_im = _RAND_2234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2235 = {1{`RANDOM}};
  _T_1297_re = _RAND_2235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2236 = {1{`RANDOM}};
  _T_1297_im = _RAND_2236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2237 = {1{`RANDOM}};
  _T_1298_re = _RAND_2237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2238 = {1{`RANDOM}};
  _T_1298_im = _RAND_2238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2239 = {1{`RANDOM}};
  _T_1299_re = _RAND_2239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2240 = {1{`RANDOM}};
  _T_1299_im = _RAND_2240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2241 = {1{`RANDOM}};
  _T_1300_re = _RAND_2241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2242 = {1{`RANDOM}};
  _T_1300_im = _RAND_2242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2243 = {1{`RANDOM}};
  _T_1301_re = _RAND_2243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2244 = {1{`RANDOM}};
  _T_1301_im = _RAND_2244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2245 = {1{`RANDOM}};
  _T_1302_re = _RAND_2245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2246 = {1{`RANDOM}};
  _T_1302_im = _RAND_2246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2247 = {1{`RANDOM}};
  _T_1303_re = _RAND_2247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2248 = {1{`RANDOM}};
  _T_1303_im = _RAND_2248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2249 = {1{`RANDOM}};
  _T_1304_re = _RAND_2249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2250 = {1{`RANDOM}};
  _T_1304_im = _RAND_2250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2251 = {1{`RANDOM}};
  _T_1305_re = _RAND_2251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2252 = {1{`RANDOM}};
  _T_1305_im = _RAND_2252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2253 = {1{`RANDOM}};
  _T_1306_re = _RAND_2253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2254 = {1{`RANDOM}};
  _T_1306_im = _RAND_2254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2255 = {1{`RANDOM}};
  _T_1307_re = _RAND_2255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2256 = {1{`RANDOM}};
  _T_1307_im = _RAND_2256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2257 = {1{`RANDOM}};
  _T_1308_re = _RAND_2257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2258 = {1{`RANDOM}};
  _T_1308_im = _RAND_2258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2259 = {1{`RANDOM}};
  _T_1309_re = _RAND_2259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2260 = {1{`RANDOM}};
  _T_1309_im = _RAND_2260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2261 = {1{`RANDOM}};
  _T_1310_re = _RAND_2261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2262 = {1{`RANDOM}};
  _T_1310_im = _RAND_2262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2263 = {1{`RANDOM}};
  _T_1311_re = _RAND_2263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2264 = {1{`RANDOM}};
  _T_1311_im = _RAND_2264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2265 = {1{`RANDOM}};
  _T_1312_re = _RAND_2265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2266 = {1{`RANDOM}};
  _T_1312_im = _RAND_2266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2267 = {1{`RANDOM}};
  _T_1313_re = _RAND_2267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2268 = {1{`RANDOM}};
  _T_1313_im = _RAND_2268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2269 = {1{`RANDOM}};
  _T_1314_re = _RAND_2269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2270 = {1{`RANDOM}};
  _T_1314_im = _RAND_2270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2271 = {1{`RANDOM}};
  _T_1315_re = _RAND_2271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2272 = {1{`RANDOM}};
  _T_1315_im = _RAND_2272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2273 = {1{`RANDOM}};
  _T_1316_re = _RAND_2273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2274 = {1{`RANDOM}};
  _T_1316_im = _RAND_2274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2275 = {1{`RANDOM}};
  _T_1317_re = _RAND_2275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2276 = {1{`RANDOM}};
  _T_1317_im = _RAND_2276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2277 = {1{`RANDOM}};
  _T_1318_re = _RAND_2277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2278 = {1{`RANDOM}};
  _T_1318_im = _RAND_2278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2279 = {1{`RANDOM}};
  _T_1319_re = _RAND_2279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2280 = {1{`RANDOM}};
  _T_1319_im = _RAND_2280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2281 = {1{`RANDOM}};
  _T_1320_re = _RAND_2281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2282 = {1{`RANDOM}};
  _T_1320_im = _RAND_2282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2283 = {1{`RANDOM}};
  _T_1321_re = _RAND_2283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2284 = {1{`RANDOM}};
  _T_1321_im = _RAND_2284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2285 = {1{`RANDOM}};
  _T_1322_re = _RAND_2285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2286 = {1{`RANDOM}};
  _T_1322_im = _RAND_2286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2287 = {1{`RANDOM}};
  _T_1323_re = _RAND_2287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2288 = {1{`RANDOM}};
  _T_1323_im = _RAND_2288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2289 = {1{`RANDOM}};
  _T_1324_re = _RAND_2289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2290 = {1{`RANDOM}};
  _T_1324_im = _RAND_2290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2291 = {1{`RANDOM}};
  _T_1325_re = _RAND_2291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2292 = {1{`RANDOM}};
  _T_1325_im = _RAND_2292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2293 = {1{`RANDOM}};
  _T_1326_re = _RAND_2293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2294 = {1{`RANDOM}};
  _T_1326_im = _RAND_2294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2295 = {1{`RANDOM}};
  _T_1327_re = _RAND_2295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2296 = {1{`RANDOM}};
  _T_1327_im = _RAND_2296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2297 = {1{`RANDOM}};
  _T_1328_re = _RAND_2297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2298 = {1{`RANDOM}};
  _T_1328_im = _RAND_2298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2299 = {1{`RANDOM}};
  _T_1329_re = _RAND_2299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2300 = {1{`RANDOM}};
  _T_1329_im = _RAND_2300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2301 = {1{`RANDOM}};
  _T_1330_re = _RAND_2301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2302 = {1{`RANDOM}};
  _T_1330_im = _RAND_2302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2303 = {1{`RANDOM}};
  _T_1331_re = _RAND_2303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2304 = {1{`RANDOM}};
  _T_1331_im = _RAND_2304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2305 = {1{`RANDOM}};
  _T_1332_re = _RAND_2305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2306 = {1{`RANDOM}};
  _T_1332_im = _RAND_2306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2307 = {1{`RANDOM}};
  _T_1333_re = _RAND_2307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2308 = {1{`RANDOM}};
  _T_1333_im = _RAND_2308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2309 = {1{`RANDOM}};
  _T_1334_re = _RAND_2309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2310 = {1{`RANDOM}};
  _T_1334_im = _RAND_2310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2311 = {1{`RANDOM}};
  _T_1335_re = _RAND_2311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2312 = {1{`RANDOM}};
  _T_1335_im = _RAND_2312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2313 = {1{`RANDOM}};
  _T_1336_re = _RAND_2313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2314 = {1{`RANDOM}};
  _T_1336_im = _RAND_2314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2315 = {1{`RANDOM}};
  _T_1337_re = _RAND_2315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2316 = {1{`RANDOM}};
  _T_1337_im = _RAND_2316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2317 = {1{`RANDOM}};
  _T_1338_re = _RAND_2317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2318 = {1{`RANDOM}};
  _T_1338_im = _RAND_2318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2319 = {1{`RANDOM}};
  _T_1339_re = _RAND_2319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2320 = {1{`RANDOM}};
  _T_1339_im = _RAND_2320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2321 = {1{`RANDOM}};
  _T_1340_re = _RAND_2321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2322 = {1{`RANDOM}};
  _T_1340_im = _RAND_2322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2323 = {1{`RANDOM}};
  _T_1341_re = _RAND_2323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2324 = {1{`RANDOM}};
  _T_1341_im = _RAND_2324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2325 = {1{`RANDOM}};
  _T_1342_re = _RAND_2325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2326 = {1{`RANDOM}};
  _T_1342_im = _RAND_2326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2327 = {1{`RANDOM}};
  _T_1343_re = _RAND_2327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2328 = {1{`RANDOM}};
  _T_1343_im = _RAND_2328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2329 = {1{`RANDOM}};
  _T_1344_re = _RAND_2329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2330 = {1{`RANDOM}};
  _T_1344_im = _RAND_2330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2331 = {1{`RANDOM}};
  _T_1345_re = _RAND_2331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2332 = {1{`RANDOM}};
  _T_1345_im = _RAND_2332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2333 = {1{`RANDOM}};
  _T_1346_re = _RAND_2333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2334 = {1{`RANDOM}};
  _T_1346_im = _RAND_2334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2335 = {1{`RANDOM}};
  _T_1347_re = _RAND_2335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2336 = {1{`RANDOM}};
  _T_1347_im = _RAND_2336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2337 = {1{`RANDOM}};
  _T_1348_re = _RAND_2337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2338 = {1{`RANDOM}};
  _T_1348_im = _RAND_2338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2339 = {1{`RANDOM}};
  _T_1349_re = _RAND_2339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2340 = {1{`RANDOM}};
  _T_1349_im = _RAND_2340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2341 = {1{`RANDOM}};
  _T_1350_re = _RAND_2341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2342 = {1{`RANDOM}};
  _T_1350_im = _RAND_2342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2343 = {1{`RANDOM}};
  _T_1351_re = _RAND_2343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2344 = {1{`RANDOM}};
  _T_1351_im = _RAND_2344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2345 = {1{`RANDOM}};
  _T_1352_re = _RAND_2345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2346 = {1{`RANDOM}};
  _T_1352_im = _RAND_2346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2347 = {1{`RANDOM}};
  _T_1353_re = _RAND_2347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2348 = {1{`RANDOM}};
  _T_1353_im = _RAND_2348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2349 = {1{`RANDOM}};
  _T_1354_re = _RAND_2349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2350 = {1{`RANDOM}};
  _T_1354_im = _RAND_2350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2351 = {1{`RANDOM}};
  _T_1355_re = _RAND_2351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2352 = {1{`RANDOM}};
  _T_1355_im = _RAND_2352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2353 = {1{`RANDOM}};
  _T_1356_re = _RAND_2353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2354 = {1{`RANDOM}};
  _T_1356_im = _RAND_2354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2355 = {1{`RANDOM}};
  _T_1357_re = _RAND_2355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2356 = {1{`RANDOM}};
  _T_1357_im = _RAND_2356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2357 = {1{`RANDOM}};
  _T_1358_re = _RAND_2357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2358 = {1{`RANDOM}};
  _T_1358_im = _RAND_2358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2359 = {1{`RANDOM}};
  _T_1359_re = _RAND_2359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2360 = {1{`RANDOM}};
  _T_1359_im = _RAND_2360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2361 = {1{`RANDOM}};
  _T_1360_re = _RAND_2361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2362 = {1{`RANDOM}};
  _T_1360_im = _RAND_2362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2363 = {1{`RANDOM}};
  _T_1361_re = _RAND_2363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2364 = {1{`RANDOM}};
  _T_1361_im = _RAND_2364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2365 = {1{`RANDOM}};
  _T_1362_re = _RAND_2365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2366 = {1{`RANDOM}};
  _T_1362_im = _RAND_2366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2367 = {1{`RANDOM}};
  _T_1363_re = _RAND_2367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2368 = {1{`RANDOM}};
  _T_1363_im = _RAND_2368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2369 = {1{`RANDOM}};
  _T_1364_re = _RAND_2369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2370 = {1{`RANDOM}};
  _T_1364_im = _RAND_2370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2371 = {1{`RANDOM}};
  _T_1365_re = _RAND_2371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2372 = {1{`RANDOM}};
  _T_1365_im = _RAND_2372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2373 = {1{`RANDOM}};
  _T_1366_re = _RAND_2373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2374 = {1{`RANDOM}};
  _T_1366_im = _RAND_2374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2375 = {1{`RANDOM}};
  _T_1367_re = _RAND_2375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2376 = {1{`RANDOM}};
  _T_1367_im = _RAND_2376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2377 = {1{`RANDOM}};
  _T_1368_re = _RAND_2377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2378 = {1{`RANDOM}};
  _T_1368_im = _RAND_2378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2379 = {1{`RANDOM}};
  _T_1369_re = _RAND_2379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2380 = {1{`RANDOM}};
  _T_1369_im = _RAND_2380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2381 = {1{`RANDOM}};
  _T_1370_re = _RAND_2381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2382 = {1{`RANDOM}};
  _T_1370_im = _RAND_2382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2383 = {1{`RANDOM}};
  _T_1371_re = _RAND_2383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2384 = {1{`RANDOM}};
  _T_1371_im = _RAND_2384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2385 = {1{`RANDOM}};
  _T_1372_re = _RAND_2385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2386 = {1{`RANDOM}};
  _T_1372_im = _RAND_2386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2387 = {1{`RANDOM}};
  _T_1373_re = _RAND_2387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2388 = {1{`RANDOM}};
  _T_1373_im = _RAND_2388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2389 = {1{`RANDOM}};
  _T_1374_re = _RAND_2389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2390 = {1{`RANDOM}};
  _T_1374_im = _RAND_2390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2391 = {1{`RANDOM}};
  _T_1375_re = _RAND_2391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2392 = {1{`RANDOM}};
  _T_1375_im = _RAND_2392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2393 = {1{`RANDOM}};
  _T_1376_re = _RAND_2393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2394 = {1{`RANDOM}};
  _T_1376_im = _RAND_2394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2395 = {1{`RANDOM}};
  _T_1377_re = _RAND_2395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2396 = {1{`RANDOM}};
  _T_1377_im = _RAND_2396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2397 = {1{`RANDOM}};
  _T_1378_re = _RAND_2397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2398 = {1{`RANDOM}};
  _T_1378_im = _RAND_2398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2399 = {1{`RANDOM}};
  _T_1379_re = _RAND_2399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2400 = {1{`RANDOM}};
  _T_1379_im = _RAND_2400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2401 = {1{`RANDOM}};
  _T_1380_re = _RAND_2401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2402 = {1{`RANDOM}};
  _T_1380_im = _RAND_2402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2403 = {1{`RANDOM}};
  _T_1381_re = _RAND_2403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2404 = {1{`RANDOM}};
  _T_1381_im = _RAND_2404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2405 = {1{`RANDOM}};
  _T_1382_re = _RAND_2405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2406 = {1{`RANDOM}};
  _T_1382_im = _RAND_2406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2407 = {1{`RANDOM}};
  _T_1383_re = _RAND_2407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2408 = {1{`RANDOM}};
  _T_1383_im = _RAND_2408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2409 = {1{`RANDOM}};
  _T_1384_re = _RAND_2409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2410 = {1{`RANDOM}};
  _T_1384_im = _RAND_2410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2411 = {1{`RANDOM}};
  _T_1385_re = _RAND_2411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2412 = {1{`RANDOM}};
  _T_1385_im = _RAND_2412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2413 = {1{`RANDOM}};
  _T_1386_re = _RAND_2413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2414 = {1{`RANDOM}};
  _T_1386_im = _RAND_2414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2415 = {1{`RANDOM}};
  _T_1387_re = _RAND_2415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2416 = {1{`RANDOM}};
  _T_1387_im = _RAND_2416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2417 = {1{`RANDOM}};
  _T_1388_re = _RAND_2417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2418 = {1{`RANDOM}};
  _T_1388_im = _RAND_2418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2419 = {1{`RANDOM}};
  _T_1389_re = _RAND_2419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2420 = {1{`RANDOM}};
  _T_1389_im = _RAND_2420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2421 = {1{`RANDOM}};
  _T_1390_re = _RAND_2421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2422 = {1{`RANDOM}};
  _T_1390_im = _RAND_2422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2423 = {1{`RANDOM}};
  _T_1391_re = _RAND_2423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2424 = {1{`RANDOM}};
  _T_1391_im = _RAND_2424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2425 = {1{`RANDOM}};
  _T_1392_re = _RAND_2425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2426 = {1{`RANDOM}};
  _T_1392_im = _RAND_2426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2427 = {1{`RANDOM}};
  _T_1393_re = _RAND_2427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2428 = {1{`RANDOM}};
  _T_1393_im = _RAND_2428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2429 = {1{`RANDOM}};
  _T_1394_re = _RAND_2429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2430 = {1{`RANDOM}};
  _T_1394_im = _RAND_2430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2431 = {1{`RANDOM}};
  _T_1395_re = _RAND_2431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2432 = {1{`RANDOM}};
  _T_1395_im = _RAND_2432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2433 = {1{`RANDOM}};
  _T_1396_re = _RAND_2433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2434 = {1{`RANDOM}};
  _T_1396_im = _RAND_2434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2435 = {1{`RANDOM}};
  _T_1397_re = _RAND_2435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2436 = {1{`RANDOM}};
  _T_1397_im = _RAND_2436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2437 = {1{`RANDOM}};
  _T_1398_re = _RAND_2437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2438 = {1{`RANDOM}};
  _T_1398_im = _RAND_2438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2439 = {1{`RANDOM}};
  _T_1399_re = _RAND_2439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2440 = {1{`RANDOM}};
  _T_1399_im = _RAND_2440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2441 = {1{`RANDOM}};
  _T_1400_re = _RAND_2441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2442 = {1{`RANDOM}};
  _T_1400_im = _RAND_2442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2443 = {1{`RANDOM}};
  _T_1401_re = _RAND_2443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2444 = {1{`RANDOM}};
  _T_1401_im = _RAND_2444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2445 = {1{`RANDOM}};
  _T_1402_re = _RAND_2445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2446 = {1{`RANDOM}};
  _T_1402_im = _RAND_2446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2447 = {1{`RANDOM}};
  _T_1403_re = _RAND_2447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2448 = {1{`RANDOM}};
  _T_1403_im = _RAND_2448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2449 = {1{`RANDOM}};
  _T_1404_re = _RAND_2449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2450 = {1{`RANDOM}};
  _T_1404_im = _RAND_2450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2451 = {1{`RANDOM}};
  _T_1405_re = _RAND_2451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2452 = {1{`RANDOM}};
  _T_1405_im = _RAND_2452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2453 = {1{`RANDOM}};
  _T_1406_re = _RAND_2453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2454 = {1{`RANDOM}};
  _T_1406_im = _RAND_2454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2455 = {1{`RANDOM}};
  _T_1407_re = _RAND_2455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2456 = {1{`RANDOM}};
  _T_1407_im = _RAND_2456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2457 = {1{`RANDOM}};
  _T_1408_re = _RAND_2457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2458 = {1{`RANDOM}};
  _T_1408_im = _RAND_2458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2459 = {1{`RANDOM}};
  _T_1409_re = _RAND_2459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2460 = {1{`RANDOM}};
  _T_1409_im = _RAND_2460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2461 = {1{`RANDOM}};
  _T_1410_re = _RAND_2461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2462 = {1{`RANDOM}};
  _T_1410_im = _RAND_2462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2463 = {1{`RANDOM}};
  _T_1411_re = _RAND_2463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2464 = {1{`RANDOM}};
  _T_1411_im = _RAND_2464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2465 = {1{`RANDOM}};
  _T_1412_re = _RAND_2465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2466 = {1{`RANDOM}};
  _T_1412_im = _RAND_2466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2467 = {1{`RANDOM}};
  _T_1413_re = _RAND_2467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2468 = {1{`RANDOM}};
  _T_1413_im = _RAND_2468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2469 = {1{`RANDOM}};
  _T_1414_re = _RAND_2469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2470 = {1{`RANDOM}};
  _T_1414_im = _RAND_2470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2471 = {1{`RANDOM}};
  _T_1415_re = _RAND_2471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2472 = {1{`RANDOM}};
  _T_1415_im = _RAND_2472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2473 = {1{`RANDOM}};
  _T_1416_re = _RAND_2473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2474 = {1{`RANDOM}};
  _T_1416_im = _RAND_2474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2475 = {1{`RANDOM}};
  _T_1417_re = _RAND_2475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2476 = {1{`RANDOM}};
  _T_1417_im = _RAND_2476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2477 = {1{`RANDOM}};
  _T_1418_re = _RAND_2477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2478 = {1{`RANDOM}};
  _T_1418_im = _RAND_2478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2479 = {1{`RANDOM}};
  _T_1419_re = _RAND_2479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2480 = {1{`RANDOM}};
  _T_1419_im = _RAND_2480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2481 = {1{`RANDOM}};
  _T_1420_re = _RAND_2481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2482 = {1{`RANDOM}};
  _T_1420_im = _RAND_2482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2483 = {1{`RANDOM}};
  _T_1421_re = _RAND_2483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2484 = {1{`RANDOM}};
  _T_1421_im = _RAND_2484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2485 = {1{`RANDOM}};
  _T_1422_re = _RAND_2485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2486 = {1{`RANDOM}};
  _T_1422_im = _RAND_2486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2487 = {1{`RANDOM}};
  _T_1423_re = _RAND_2487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2488 = {1{`RANDOM}};
  _T_1423_im = _RAND_2488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2489 = {1{`RANDOM}};
  _T_1424_re = _RAND_2489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2490 = {1{`RANDOM}};
  _T_1424_im = _RAND_2490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2491 = {1{`RANDOM}};
  _T_1425_re = _RAND_2491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2492 = {1{`RANDOM}};
  _T_1425_im = _RAND_2492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2493 = {1{`RANDOM}};
  _T_1426_re = _RAND_2493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2494 = {1{`RANDOM}};
  _T_1426_im = _RAND_2494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2495 = {1{`RANDOM}};
  _T_1427_re = _RAND_2495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2496 = {1{`RANDOM}};
  _T_1427_im = _RAND_2496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2497 = {1{`RANDOM}};
  _T_1428_re = _RAND_2497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2498 = {1{`RANDOM}};
  _T_1428_im = _RAND_2498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2499 = {1{`RANDOM}};
  _T_1429_re = _RAND_2499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2500 = {1{`RANDOM}};
  _T_1429_im = _RAND_2500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2501 = {1{`RANDOM}};
  _T_1430_re = _RAND_2501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2502 = {1{`RANDOM}};
  _T_1430_im = _RAND_2502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2503 = {1{`RANDOM}};
  _T_1431_re = _RAND_2503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2504 = {1{`RANDOM}};
  _T_1431_im = _RAND_2504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2505 = {1{`RANDOM}};
  _T_1432_re = _RAND_2505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2506 = {1{`RANDOM}};
  _T_1432_im = _RAND_2506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2507 = {1{`RANDOM}};
  _T_1433_re = _RAND_2507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2508 = {1{`RANDOM}};
  _T_1433_im = _RAND_2508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2509 = {1{`RANDOM}};
  _T_1434_re = _RAND_2509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2510 = {1{`RANDOM}};
  _T_1434_im = _RAND_2510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2511 = {1{`RANDOM}};
  _T_1435_re = _RAND_2511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2512 = {1{`RANDOM}};
  _T_1435_im = _RAND_2512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2513 = {1{`RANDOM}};
  _T_1436_re = _RAND_2513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2514 = {1{`RANDOM}};
  _T_1436_im = _RAND_2514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2515 = {1{`RANDOM}};
  _T_1437_re = _RAND_2515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2516 = {1{`RANDOM}};
  _T_1437_im = _RAND_2516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2517 = {1{`RANDOM}};
  _T_1438_re = _RAND_2517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2518 = {1{`RANDOM}};
  _T_1438_im = _RAND_2518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2519 = {1{`RANDOM}};
  _T_1439_re = _RAND_2519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2520 = {1{`RANDOM}};
  _T_1439_im = _RAND_2520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2521 = {1{`RANDOM}};
  _T_1440_re = _RAND_2521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2522 = {1{`RANDOM}};
  _T_1440_im = _RAND_2522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2523 = {1{`RANDOM}};
  _T_1441_re = _RAND_2523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2524 = {1{`RANDOM}};
  _T_1441_im = _RAND_2524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2525 = {1{`RANDOM}};
  _T_1442_re = _RAND_2525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2526 = {1{`RANDOM}};
  _T_1442_im = _RAND_2526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2527 = {1{`RANDOM}};
  _T_1443_re = _RAND_2527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2528 = {1{`RANDOM}};
  _T_1443_im = _RAND_2528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2529 = {1{`RANDOM}};
  _T_1444_re = _RAND_2529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2530 = {1{`RANDOM}};
  _T_1444_im = _RAND_2530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2531 = {1{`RANDOM}};
  _T_1445_re = _RAND_2531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2532 = {1{`RANDOM}};
  _T_1445_im = _RAND_2532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2533 = {1{`RANDOM}};
  _T_1446_re = _RAND_2533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2534 = {1{`RANDOM}};
  _T_1446_im = _RAND_2534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2535 = {1{`RANDOM}};
  _T_1447_re = _RAND_2535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2536 = {1{`RANDOM}};
  _T_1447_im = _RAND_2536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2537 = {1{`RANDOM}};
  _T_1448_re = _RAND_2537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2538 = {1{`RANDOM}};
  _T_1448_im = _RAND_2538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2539 = {1{`RANDOM}};
  _T_1449_re = _RAND_2539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2540 = {1{`RANDOM}};
  _T_1449_im = _RAND_2540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2541 = {1{`RANDOM}};
  _T_1450_re = _RAND_2541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2542 = {1{`RANDOM}};
  _T_1450_im = _RAND_2542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2543 = {1{`RANDOM}};
  _T_1451_re = _RAND_2543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2544 = {1{`RANDOM}};
  _T_1451_im = _RAND_2544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2545 = {1{`RANDOM}};
  _T_1452_re = _RAND_2545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2546 = {1{`RANDOM}};
  _T_1452_im = _RAND_2546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2547 = {1{`RANDOM}};
  _T_1453_re = _RAND_2547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2548 = {1{`RANDOM}};
  _T_1453_im = _RAND_2548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2549 = {1{`RANDOM}};
  _T_1454_re = _RAND_2549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2550 = {1{`RANDOM}};
  _T_1454_im = _RAND_2550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2551 = {1{`RANDOM}};
  _T_1455_re = _RAND_2551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2552 = {1{`RANDOM}};
  _T_1455_im = _RAND_2552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2553 = {1{`RANDOM}};
  _T_1456_re = _RAND_2553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2554 = {1{`RANDOM}};
  _T_1456_im = _RAND_2554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2555 = {1{`RANDOM}};
  _T_1457_re = _RAND_2555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2556 = {1{`RANDOM}};
  _T_1457_im = _RAND_2556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2557 = {1{`RANDOM}};
  _T_1458_re = _RAND_2557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2558 = {1{`RANDOM}};
  _T_1458_im = _RAND_2558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2559 = {1{`RANDOM}};
  _T_1459_re = _RAND_2559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2560 = {1{`RANDOM}};
  _T_1459_im = _RAND_2560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2561 = {1{`RANDOM}};
  _T_1460_re = _RAND_2561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2562 = {1{`RANDOM}};
  _T_1460_im = _RAND_2562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2563 = {1{`RANDOM}};
  _T_1461_re = _RAND_2563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2564 = {1{`RANDOM}};
  _T_1461_im = _RAND_2564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2565 = {1{`RANDOM}};
  _T_1462_re = _RAND_2565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2566 = {1{`RANDOM}};
  _T_1462_im = _RAND_2566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2567 = {1{`RANDOM}};
  _T_1463_re = _RAND_2567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2568 = {1{`RANDOM}};
  _T_1463_im = _RAND_2568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2569 = {1{`RANDOM}};
  _T_1464_re = _RAND_2569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2570 = {1{`RANDOM}};
  _T_1464_im = _RAND_2570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2571 = {1{`RANDOM}};
  _T_1465_re = _RAND_2571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2572 = {1{`RANDOM}};
  _T_1465_im = _RAND_2572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2573 = {1{`RANDOM}};
  _T_1466_re = _RAND_2573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2574 = {1{`RANDOM}};
  _T_1466_im = _RAND_2574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2575 = {1{`RANDOM}};
  _T_1467_re = _RAND_2575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2576 = {1{`RANDOM}};
  _T_1467_im = _RAND_2576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2577 = {1{`RANDOM}};
  _T_1468_re = _RAND_2577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2578 = {1{`RANDOM}};
  _T_1468_im = _RAND_2578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2579 = {1{`RANDOM}};
  _T_1469_re = _RAND_2579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2580 = {1{`RANDOM}};
  _T_1469_im = _RAND_2580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2581 = {1{`RANDOM}};
  _T_1470_re = _RAND_2581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2582 = {1{`RANDOM}};
  _T_1470_im = _RAND_2582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2583 = {1{`RANDOM}};
  _T_1471_re = _RAND_2583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2584 = {1{`RANDOM}};
  _T_1471_im = _RAND_2584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2585 = {1{`RANDOM}};
  _T_1472_re = _RAND_2585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2586 = {1{`RANDOM}};
  _T_1472_im = _RAND_2586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2587 = {1{`RANDOM}};
  _T_1473_re = _RAND_2587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2588 = {1{`RANDOM}};
  _T_1473_im = _RAND_2588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2589 = {1{`RANDOM}};
  _T_1474_re = _RAND_2589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2590 = {1{`RANDOM}};
  _T_1474_im = _RAND_2590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2591 = {1{`RANDOM}};
  _T_1475_re = _RAND_2591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2592 = {1{`RANDOM}};
  _T_1475_im = _RAND_2592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2593 = {1{`RANDOM}};
  _T_1476_re = _RAND_2593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2594 = {1{`RANDOM}};
  _T_1476_im = _RAND_2594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2595 = {1{`RANDOM}};
  _T_1477_re = _RAND_2595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2596 = {1{`RANDOM}};
  _T_1477_im = _RAND_2596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2597 = {1{`RANDOM}};
  _T_1478_re = _RAND_2597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2598 = {1{`RANDOM}};
  _T_1478_im = _RAND_2598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2599 = {1{`RANDOM}};
  _T_1479_re = _RAND_2599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2600 = {1{`RANDOM}};
  _T_1479_im = _RAND_2600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2601 = {1{`RANDOM}};
  _T_1480_re = _RAND_2601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2602 = {1{`RANDOM}};
  _T_1480_im = _RAND_2602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2603 = {1{`RANDOM}};
  _T_1481_re = _RAND_2603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2604 = {1{`RANDOM}};
  _T_1481_im = _RAND_2604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2605 = {1{`RANDOM}};
  _T_1482_re = _RAND_2605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2606 = {1{`RANDOM}};
  _T_1482_im = _RAND_2606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2607 = {1{`RANDOM}};
  _T_1483_re = _RAND_2607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2608 = {1{`RANDOM}};
  _T_1483_im = _RAND_2608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2609 = {1{`RANDOM}};
  _T_1484_re = _RAND_2609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2610 = {1{`RANDOM}};
  _T_1484_im = _RAND_2610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2611 = {1{`RANDOM}};
  _T_1485_re = _RAND_2611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2612 = {1{`RANDOM}};
  _T_1485_im = _RAND_2612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2613 = {1{`RANDOM}};
  _T_1486_re = _RAND_2613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2614 = {1{`RANDOM}};
  _T_1486_im = _RAND_2614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2615 = {1{`RANDOM}};
  _T_1487_re = _RAND_2615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2616 = {1{`RANDOM}};
  _T_1487_im = _RAND_2616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2617 = {1{`RANDOM}};
  _T_1488_re = _RAND_2617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2618 = {1{`RANDOM}};
  _T_1488_im = _RAND_2618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2619 = {1{`RANDOM}};
  _T_1489_re = _RAND_2619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2620 = {1{`RANDOM}};
  _T_1489_im = _RAND_2620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2621 = {1{`RANDOM}};
  _T_1490_re = _RAND_2621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2622 = {1{`RANDOM}};
  _T_1490_im = _RAND_2622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2623 = {1{`RANDOM}};
  _T_1491_re = _RAND_2623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2624 = {1{`RANDOM}};
  _T_1491_im = _RAND_2624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2625 = {1{`RANDOM}};
  _T_1492_re = _RAND_2625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2626 = {1{`RANDOM}};
  _T_1492_im = _RAND_2626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2627 = {1{`RANDOM}};
  _T_1493_re = _RAND_2627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2628 = {1{`RANDOM}};
  _T_1493_im = _RAND_2628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2629 = {1{`RANDOM}};
  _T_1494_re = _RAND_2629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2630 = {1{`RANDOM}};
  _T_1494_im = _RAND_2630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2631 = {1{`RANDOM}};
  _T_1495_re = _RAND_2631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2632 = {1{`RANDOM}};
  _T_1495_im = _RAND_2632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2633 = {1{`RANDOM}};
  _T_1496_re = _RAND_2633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2634 = {1{`RANDOM}};
  _T_1496_im = _RAND_2634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2635 = {1{`RANDOM}};
  _T_1497_re = _RAND_2635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2636 = {1{`RANDOM}};
  _T_1497_im = _RAND_2636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2637 = {1{`RANDOM}};
  _T_1498_re = _RAND_2637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2638 = {1{`RANDOM}};
  _T_1498_im = _RAND_2638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2639 = {1{`RANDOM}};
  _T_1499_re = _RAND_2639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2640 = {1{`RANDOM}};
  _T_1499_im = _RAND_2640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2641 = {1{`RANDOM}};
  _T_1500_re = _RAND_2641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2642 = {1{`RANDOM}};
  _T_1500_im = _RAND_2642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2643 = {1{`RANDOM}};
  _T_1501_re = _RAND_2643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2644 = {1{`RANDOM}};
  _T_1501_im = _RAND_2644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2645 = {1{`RANDOM}};
  _T_1502_re = _RAND_2645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2646 = {1{`RANDOM}};
  _T_1502_im = _RAND_2646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2647 = {1{`RANDOM}};
  _T_1503_re = _RAND_2647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2648 = {1{`RANDOM}};
  _T_1503_im = _RAND_2648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2649 = {1{`RANDOM}};
  _T_1504_re = _RAND_2649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2650 = {1{`RANDOM}};
  _T_1504_im = _RAND_2650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2651 = {1{`RANDOM}};
  _T_1505_re = _RAND_2651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2652 = {1{`RANDOM}};
  _T_1505_im = _RAND_2652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2653 = {1{`RANDOM}};
  _T_1506_re = _RAND_2653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2654 = {1{`RANDOM}};
  _T_1506_im = _RAND_2654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2655 = {1{`RANDOM}};
  _T_1507_re = _RAND_2655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2656 = {1{`RANDOM}};
  _T_1507_im = _RAND_2656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2657 = {1{`RANDOM}};
  _T_1508_re = _RAND_2657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2658 = {1{`RANDOM}};
  _T_1508_im = _RAND_2658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2659 = {1{`RANDOM}};
  _T_1509_re = _RAND_2659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2660 = {1{`RANDOM}};
  _T_1509_im = _RAND_2660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2661 = {1{`RANDOM}};
  _T_1510_re = _RAND_2661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2662 = {1{`RANDOM}};
  _T_1510_im = _RAND_2662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2663 = {1{`RANDOM}};
  _T_1511_re = _RAND_2663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2664 = {1{`RANDOM}};
  _T_1511_im = _RAND_2664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2665 = {1{`RANDOM}};
  _T_1512_re = _RAND_2665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2666 = {1{`RANDOM}};
  _T_1512_im = _RAND_2666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2667 = {1{`RANDOM}};
  _T_1513_re = _RAND_2667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2668 = {1{`RANDOM}};
  _T_1513_im = _RAND_2668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2669 = {1{`RANDOM}};
  _T_1514_re = _RAND_2669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2670 = {1{`RANDOM}};
  _T_1514_im = _RAND_2670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2671 = {1{`RANDOM}};
  _T_1515_re = _RAND_2671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2672 = {1{`RANDOM}};
  _T_1515_im = _RAND_2672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2673 = {1{`RANDOM}};
  _T_1516_re = _RAND_2673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2674 = {1{`RANDOM}};
  _T_1516_im = _RAND_2674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2675 = {1{`RANDOM}};
  _T_1517_re = _RAND_2675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2676 = {1{`RANDOM}};
  _T_1517_im = _RAND_2676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2677 = {1{`RANDOM}};
  _T_1518_re = _RAND_2677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2678 = {1{`RANDOM}};
  _T_1518_im = _RAND_2678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2679 = {1{`RANDOM}};
  _T_1519_re = _RAND_2679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2680 = {1{`RANDOM}};
  _T_1519_im = _RAND_2680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2681 = {1{`RANDOM}};
  _T_1520_re = _RAND_2681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2682 = {1{`RANDOM}};
  _T_1520_im = _RAND_2682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2683 = {1{`RANDOM}};
  _T_1521_re = _RAND_2683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2684 = {1{`RANDOM}};
  _T_1521_im = _RAND_2684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2685 = {1{`RANDOM}};
  _T_1522_re = _RAND_2685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2686 = {1{`RANDOM}};
  _T_1522_im = _RAND_2686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2687 = {1{`RANDOM}};
  _T_1523_re = _RAND_2687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2688 = {1{`RANDOM}};
  _T_1523_im = _RAND_2688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2689 = {1{`RANDOM}};
  _T_1524_re = _RAND_2689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2690 = {1{`RANDOM}};
  _T_1524_im = _RAND_2690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2691 = {1{`RANDOM}};
  _T_1525_re = _RAND_2691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2692 = {1{`RANDOM}};
  _T_1525_im = _RAND_2692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2693 = {1{`RANDOM}};
  _T_1526_re = _RAND_2693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2694 = {1{`RANDOM}};
  _T_1526_im = _RAND_2694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2695 = {1{`RANDOM}};
  _T_1527_re = _RAND_2695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2696 = {1{`RANDOM}};
  _T_1527_im = _RAND_2696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2697 = {1{`RANDOM}};
  _T_1528_re = _RAND_2697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2698 = {1{`RANDOM}};
  _T_1528_im = _RAND_2698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2699 = {1{`RANDOM}};
  _T_1529_re = _RAND_2699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2700 = {1{`RANDOM}};
  _T_1529_im = _RAND_2700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2701 = {1{`RANDOM}};
  _T_1530_re = _RAND_2701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2702 = {1{`RANDOM}};
  _T_1530_im = _RAND_2702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2703 = {1{`RANDOM}};
  _T_1531_re = _RAND_2703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2704 = {1{`RANDOM}};
  _T_1531_im = _RAND_2704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2705 = {1{`RANDOM}};
  _T_1532_re = _RAND_2705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2706 = {1{`RANDOM}};
  _T_1532_im = _RAND_2706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2707 = {1{`RANDOM}};
  _T_1533_re = _RAND_2707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2708 = {1{`RANDOM}};
  _T_1533_im = _RAND_2708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2709 = {1{`RANDOM}};
  _T_1534_re = _RAND_2709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2710 = {1{`RANDOM}};
  _T_1534_im = _RAND_2710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2711 = {1{`RANDOM}};
  _T_1535_re = _RAND_2711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2712 = {1{`RANDOM}};
  _T_1535_im = _RAND_2712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2713 = {1{`RANDOM}};
  _T_1536_re = _RAND_2713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2714 = {1{`RANDOM}};
  _T_1536_im = _RAND_2714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2715 = {1{`RANDOM}};
  _T_1537_re = _RAND_2715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2716 = {1{`RANDOM}};
  _T_1537_im = _RAND_2716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2717 = {1{`RANDOM}};
  _T_1538_re = _RAND_2717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2718 = {1{`RANDOM}};
  _T_1538_im = _RAND_2718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2719 = {1{`RANDOM}};
  _T_1539_re = _RAND_2719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2720 = {1{`RANDOM}};
  _T_1539_im = _RAND_2720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2721 = {1{`RANDOM}};
  _T_1540_re = _RAND_2721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2722 = {1{`RANDOM}};
  _T_1540_im = _RAND_2722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2723 = {1{`RANDOM}};
  _T_1541_re = _RAND_2723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2724 = {1{`RANDOM}};
  _T_1541_im = _RAND_2724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2725 = {1{`RANDOM}};
  _T_1542_re = _RAND_2725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2726 = {1{`RANDOM}};
  _T_1542_im = _RAND_2726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2727 = {1{`RANDOM}};
  _T_1543_re = _RAND_2727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2728 = {1{`RANDOM}};
  _T_1543_im = _RAND_2728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2729 = {1{`RANDOM}};
  _T_1544_re = _RAND_2729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2730 = {1{`RANDOM}};
  _T_1544_im = _RAND_2730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2731 = {1{`RANDOM}};
  _T_1545_re = _RAND_2731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2732 = {1{`RANDOM}};
  _T_1545_im = _RAND_2732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2733 = {1{`RANDOM}};
  _T_1546_re = _RAND_2733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2734 = {1{`RANDOM}};
  _T_1546_im = _RAND_2734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2735 = {1{`RANDOM}};
  _T_1547_re = _RAND_2735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2736 = {1{`RANDOM}};
  _T_1547_im = _RAND_2736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2737 = {1{`RANDOM}};
  _T_1548_re = _RAND_2737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2738 = {1{`RANDOM}};
  _T_1548_im = _RAND_2738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2739 = {1{`RANDOM}};
  _T_1549_re = _RAND_2739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2740 = {1{`RANDOM}};
  _T_1549_im = _RAND_2740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2741 = {1{`RANDOM}};
  _T_1550_re = _RAND_2741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2742 = {1{`RANDOM}};
  _T_1550_im = _RAND_2742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2743 = {1{`RANDOM}};
  _T_1551_re = _RAND_2743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2744 = {1{`RANDOM}};
  _T_1551_im = _RAND_2744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2745 = {1{`RANDOM}};
  _T_1552_re = _RAND_2745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2746 = {1{`RANDOM}};
  _T_1552_im = _RAND_2746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2747 = {1{`RANDOM}};
  _T_1553_re = _RAND_2747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2748 = {1{`RANDOM}};
  _T_1553_im = _RAND_2748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2749 = {1{`RANDOM}};
  _T_1554_re = _RAND_2749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2750 = {1{`RANDOM}};
  _T_1554_im = _RAND_2750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2751 = {1{`RANDOM}};
  _T_1555_re = _RAND_2751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2752 = {1{`RANDOM}};
  _T_1555_im = _RAND_2752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2753 = {1{`RANDOM}};
  _T_1556_re = _RAND_2753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2754 = {1{`RANDOM}};
  _T_1556_im = _RAND_2754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2755 = {1{`RANDOM}};
  _T_1557_re = _RAND_2755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2756 = {1{`RANDOM}};
  _T_1557_im = _RAND_2756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2757 = {1{`RANDOM}};
  _T_1558_re = _RAND_2757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2758 = {1{`RANDOM}};
  _T_1558_im = _RAND_2758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2759 = {1{`RANDOM}};
  _T_1559_re = _RAND_2759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2760 = {1{`RANDOM}};
  _T_1559_im = _RAND_2760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2761 = {1{`RANDOM}};
  _T_1560_re = _RAND_2761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2762 = {1{`RANDOM}};
  _T_1560_im = _RAND_2762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2763 = {1{`RANDOM}};
  _T_1561_re = _RAND_2763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2764 = {1{`RANDOM}};
  _T_1561_im = _RAND_2764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2765 = {1{`RANDOM}};
  _T_1562_re = _RAND_2765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2766 = {1{`RANDOM}};
  _T_1562_im = _RAND_2766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2767 = {1{`RANDOM}};
  _T_1563_re = _RAND_2767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2768 = {1{`RANDOM}};
  _T_1563_im = _RAND_2768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2769 = {1{`RANDOM}};
  _T_1564_re = _RAND_2769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2770 = {1{`RANDOM}};
  _T_1564_im = _RAND_2770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2771 = {1{`RANDOM}};
  _T_1565_re = _RAND_2771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2772 = {1{`RANDOM}};
  _T_1565_im = _RAND_2772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2773 = {1{`RANDOM}};
  _T_1566_re = _RAND_2773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2774 = {1{`RANDOM}};
  _T_1566_im = _RAND_2774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2775 = {1{`RANDOM}};
  _T_1567_re = _RAND_2775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2776 = {1{`RANDOM}};
  _T_1567_im = _RAND_2776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2777 = {1{`RANDOM}};
  _T_1568_re = _RAND_2777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2778 = {1{`RANDOM}};
  _T_1568_im = _RAND_2778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2779 = {1{`RANDOM}};
  _T_1569_re = _RAND_2779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2780 = {1{`RANDOM}};
  _T_1569_im = _RAND_2780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2781 = {1{`RANDOM}};
  _T_1570_re = _RAND_2781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2782 = {1{`RANDOM}};
  _T_1570_im = _RAND_2782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2783 = {1{`RANDOM}};
  _T_1571_re = _RAND_2783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2784 = {1{`RANDOM}};
  _T_1571_im = _RAND_2784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2785 = {1{`RANDOM}};
  _T_1572_re = _RAND_2785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2786 = {1{`RANDOM}};
  _T_1572_im = _RAND_2786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2787 = {1{`RANDOM}};
  _T_1573_re = _RAND_2787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2788 = {1{`RANDOM}};
  _T_1573_im = _RAND_2788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2789 = {1{`RANDOM}};
  _T_1574_re = _RAND_2789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2790 = {1{`RANDOM}};
  _T_1574_im = _RAND_2790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2791 = {1{`RANDOM}};
  _T_1575_re = _RAND_2791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2792 = {1{`RANDOM}};
  _T_1575_im = _RAND_2792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2793 = {1{`RANDOM}};
  _T_1576_re = _RAND_2793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2794 = {1{`RANDOM}};
  _T_1576_im = _RAND_2794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2795 = {1{`RANDOM}};
  _T_1577_re = _RAND_2795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2796 = {1{`RANDOM}};
  _T_1577_im = _RAND_2796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2797 = {1{`RANDOM}};
  _T_1578_re = _RAND_2797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2798 = {1{`RANDOM}};
  _T_1578_im = _RAND_2798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2799 = {1{`RANDOM}};
  _T_1579_re = _RAND_2799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2800 = {1{`RANDOM}};
  _T_1579_im = _RAND_2800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2801 = {1{`RANDOM}};
  _T_1580_re = _RAND_2801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2802 = {1{`RANDOM}};
  _T_1580_im = _RAND_2802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2803 = {1{`RANDOM}};
  _T_1581_re = _RAND_2803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2804 = {1{`RANDOM}};
  _T_1581_im = _RAND_2804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2805 = {1{`RANDOM}};
  _T_1582_re = _RAND_2805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2806 = {1{`RANDOM}};
  _T_1582_im = _RAND_2806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2807 = {1{`RANDOM}};
  _T_1583_re = _RAND_2807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2808 = {1{`RANDOM}};
  _T_1583_im = _RAND_2808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2809 = {1{`RANDOM}};
  _T_1584_re = _RAND_2809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2810 = {1{`RANDOM}};
  _T_1584_im = _RAND_2810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2811 = {1{`RANDOM}};
  _T_1585_re = _RAND_2811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2812 = {1{`RANDOM}};
  _T_1585_im = _RAND_2812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2813 = {1{`RANDOM}};
  _T_1586_re = _RAND_2813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2814 = {1{`RANDOM}};
  _T_1586_im = _RAND_2814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2815 = {1{`RANDOM}};
  _T_1587_re = _RAND_2815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2816 = {1{`RANDOM}};
  _T_1587_im = _RAND_2816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2817 = {1{`RANDOM}};
  _T_1588_re = _RAND_2817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2818 = {1{`RANDOM}};
  _T_1588_im = _RAND_2818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2819 = {1{`RANDOM}};
  _T_1589_re = _RAND_2819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2820 = {1{`RANDOM}};
  _T_1589_im = _RAND_2820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2821 = {1{`RANDOM}};
  _T_1590_re = _RAND_2821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2822 = {1{`RANDOM}};
  _T_1590_im = _RAND_2822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2823 = {1{`RANDOM}};
  _T_1591_re = _RAND_2823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2824 = {1{`RANDOM}};
  _T_1591_im = _RAND_2824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2825 = {1{`RANDOM}};
  _T_1592_re = _RAND_2825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2826 = {1{`RANDOM}};
  _T_1592_im = _RAND_2826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2827 = {1{`RANDOM}};
  _T_1593_re = _RAND_2827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2828 = {1{`RANDOM}};
  _T_1593_im = _RAND_2828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2829 = {1{`RANDOM}};
  _T_1594_re = _RAND_2829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2830 = {1{`RANDOM}};
  _T_1594_im = _RAND_2830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2831 = {1{`RANDOM}};
  _T_1595_re = _RAND_2831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2832 = {1{`RANDOM}};
  _T_1595_im = _RAND_2832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2833 = {1{`RANDOM}};
  _T_1596_re = _RAND_2833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2834 = {1{`RANDOM}};
  _T_1596_im = _RAND_2834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2835 = {1{`RANDOM}};
  _T_1597_re = _RAND_2835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2836 = {1{`RANDOM}};
  _T_1597_im = _RAND_2836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2837 = {1{`RANDOM}};
  _T_1598_re = _RAND_2837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2838 = {1{`RANDOM}};
  _T_1598_im = _RAND_2838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2839 = {1{`RANDOM}};
  _T_1599_re = _RAND_2839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2840 = {1{`RANDOM}};
  _T_1599_im = _RAND_2840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2841 = {1{`RANDOM}};
  _T_1600_re = _RAND_2841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2842 = {1{`RANDOM}};
  _T_1600_im = _RAND_2842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2843 = {1{`RANDOM}};
  _T_1601_re = _RAND_2843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2844 = {1{`RANDOM}};
  _T_1601_im = _RAND_2844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2845 = {1{`RANDOM}};
  _T_1602_re = _RAND_2845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2846 = {1{`RANDOM}};
  _T_1602_im = _RAND_2846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2847 = {1{`RANDOM}};
  _T_1603_re = _RAND_2847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2848 = {1{`RANDOM}};
  _T_1603_im = _RAND_2848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2849 = {1{`RANDOM}};
  _T_1604_re = _RAND_2849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2850 = {1{`RANDOM}};
  _T_1604_im = _RAND_2850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2851 = {1{`RANDOM}};
  _T_1605_re = _RAND_2851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2852 = {1{`RANDOM}};
  _T_1605_im = _RAND_2852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2853 = {1{`RANDOM}};
  _T_1606_re = _RAND_2853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2854 = {1{`RANDOM}};
  _T_1606_im = _RAND_2854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2855 = {1{`RANDOM}};
  _T_1607_re = _RAND_2855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2856 = {1{`RANDOM}};
  _T_1607_im = _RAND_2856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2857 = {1{`RANDOM}};
  _T_1608_re = _RAND_2857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2858 = {1{`RANDOM}};
  _T_1608_im = _RAND_2858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2859 = {1{`RANDOM}};
  _T_1609_re = _RAND_2859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2860 = {1{`RANDOM}};
  _T_1609_im = _RAND_2860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2861 = {1{`RANDOM}};
  _T_1610_re = _RAND_2861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2862 = {1{`RANDOM}};
  _T_1610_im = _RAND_2862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2863 = {1{`RANDOM}};
  _T_1611_re = _RAND_2863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2864 = {1{`RANDOM}};
  _T_1611_im = _RAND_2864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2865 = {1{`RANDOM}};
  _T_1612_re = _RAND_2865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2866 = {1{`RANDOM}};
  _T_1612_im = _RAND_2866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2867 = {1{`RANDOM}};
  _T_1613_re = _RAND_2867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2868 = {1{`RANDOM}};
  _T_1613_im = _RAND_2868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2869 = {1{`RANDOM}};
  _T_1614_re = _RAND_2869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2870 = {1{`RANDOM}};
  _T_1614_im = _RAND_2870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2871 = {1{`RANDOM}};
  _T_1615_re = _RAND_2871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2872 = {1{`RANDOM}};
  _T_1615_im = _RAND_2872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2873 = {1{`RANDOM}};
  _T_1616_re = _RAND_2873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2874 = {1{`RANDOM}};
  _T_1616_im = _RAND_2874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2875 = {1{`RANDOM}};
  _T_1617_re = _RAND_2875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2876 = {1{`RANDOM}};
  _T_1617_im = _RAND_2876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2877 = {1{`RANDOM}};
  _T_1618_re = _RAND_2877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2878 = {1{`RANDOM}};
  _T_1618_im = _RAND_2878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2879 = {1{`RANDOM}};
  _T_1619_re = _RAND_2879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2880 = {1{`RANDOM}};
  _T_1619_im = _RAND_2880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2881 = {1{`RANDOM}};
  _T_1620_re = _RAND_2881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2882 = {1{`RANDOM}};
  _T_1620_im = _RAND_2882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2883 = {1{`RANDOM}};
  _T_1621_re = _RAND_2883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2884 = {1{`RANDOM}};
  _T_1621_im = _RAND_2884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2885 = {1{`RANDOM}};
  _T_1622_re = _RAND_2885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2886 = {1{`RANDOM}};
  _T_1622_im = _RAND_2886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2887 = {1{`RANDOM}};
  _T_1623_re = _RAND_2887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2888 = {1{`RANDOM}};
  _T_1623_im = _RAND_2888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2889 = {1{`RANDOM}};
  _T_1624_re = _RAND_2889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2890 = {1{`RANDOM}};
  _T_1624_im = _RAND_2890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2891 = {1{`RANDOM}};
  _T_1625_re = _RAND_2891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2892 = {1{`RANDOM}};
  _T_1625_im = _RAND_2892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2893 = {1{`RANDOM}};
  _T_1626_re = _RAND_2893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2894 = {1{`RANDOM}};
  _T_1626_im = _RAND_2894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2895 = {1{`RANDOM}};
  _T_1627_re = _RAND_2895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2896 = {1{`RANDOM}};
  _T_1627_im = _RAND_2896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2897 = {1{`RANDOM}};
  _T_1628_re = _RAND_2897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2898 = {1{`RANDOM}};
  _T_1628_im = _RAND_2898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2899 = {1{`RANDOM}};
  _T_1629_re = _RAND_2899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2900 = {1{`RANDOM}};
  _T_1629_im = _RAND_2900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2901 = {1{`RANDOM}};
  _T_1630_re = _RAND_2901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2902 = {1{`RANDOM}};
  _T_1630_im = _RAND_2902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2903 = {1{`RANDOM}};
  _T_1631_re = _RAND_2903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2904 = {1{`RANDOM}};
  _T_1631_im = _RAND_2904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2905 = {1{`RANDOM}};
  _T_1632_re = _RAND_2905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2906 = {1{`RANDOM}};
  _T_1632_im = _RAND_2906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2907 = {1{`RANDOM}};
  _T_1633_re = _RAND_2907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2908 = {1{`RANDOM}};
  _T_1633_im = _RAND_2908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2909 = {1{`RANDOM}};
  _T_1634_re = _RAND_2909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2910 = {1{`RANDOM}};
  _T_1634_im = _RAND_2910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2911 = {1{`RANDOM}};
  _T_1635_re = _RAND_2911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2912 = {1{`RANDOM}};
  _T_1635_im = _RAND_2912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2913 = {1{`RANDOM}};
  _T_1636_re = _RAND_2913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2914 = {1{`RANDOM}};
  _T_1636_im = _RAND_2914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2915 = {1{`RANDOM}};
  _T_1637_re = _RAND_2915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2916 = {1{`RANDOM}};
  _T_1637_im = _RAND_2916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2917 = {1{`RANDOM}};
  _T_1638_re = _RAND_2917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2918 = {1{`RANDOM}};
  _T_1638_im = _RAND_2918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2919 = {1{`RANDOM}};
  _T_1639_re = _RAND_2919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2920 = {1{`RANDOM}};
  _T_1639_im = _RAND_2920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2921 = {1{`RANDOM}};
  _T_1640_re = _RAND_2921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2922 = {1{`RANDOM}};
  _T_1640_im = _RAND_2922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2923 = {1{`RANDOM}};
  _T_1641_re = _RAND_2923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2924 = {1{`RANDOM}};
  _T_1641_im = _RAND_2924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2925 = {1{`RANDOM}};
  _T_1642_re = _RAND_2925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2926 = {1{`RANDOM}};
  _T_1642_im = _RAND_2926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2927 = {1{`RANDOM}};
  _T_1643_re = _RAND_2927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2928 = {1{`RANDOM}};
  _T_1643_im = _RAND_2928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2929 = {1{`RANDOM}};
  _T_1644_re = _RAND_2929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2930 = {1{`RANDOM}};
  _T_1644_im = _RAND_2930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2931 = {1{`RANDOM}};
  _T_1645_re = _RAND_2931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2932 = {1{`RANDOM}};
  _T_1645_im = _RAND_2932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2933 = {1{`RANDOM}};
  _T_1646_re = _RAND_2933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2934 = {1{`RANDOM}};
  _T_1646_im = _RAND_2934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2935 = {1{`RANDOM}};
  _T_1647_re = _RAND_2935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2936 = {1{`RANDOM}};
  _T_1647_im = _RAND_2936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2937 = {1{`RANDOM}};
  _T_1648_re = _RAND_2937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2938 = {1{`RANDOM}};
  _T_1648_im = _RAND_2938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2939 = {1{`RANDOM}};
  _T_1649_re = _RAND_2939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2940 = {1{`RANDOM}};
  _T_1649_im = _RAND_2940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2941 = {1{`RANDOM}};
  _T_1650_re = _RAND_2941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2942 = {1{`RANDOM}};
  _T_1650_im = _RAND_2942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2943 = {1{`RANDOM}};
  _T_1651_re = _RAND_2943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2944 = {1{`RANDOM}};
  _T_1651_im = _RAND_2944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2945 = {1{`RANDOM}};
  _T_1652_re = _RAND_2945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2946 = {1{`RANDOM}};
  _T_1652_im = _RAND_2946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2947 = {1{`RANDOM}};
  _T_1653_re = _RAND_2947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2948 = {1{`RANDOM}};
  _T_1653_im = _RAND_2948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2949 = {1{`RANDOM}};
  _T_1654_re = _RAND_2949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2950 = {1{`RANDOM}};
  _T_1654_im = _RAND_2950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2951 = {1{`RANDOM}};
  _T_1655_re = _RAND_2951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2952 = {1{`RANDOM}};
  _T_1655_im = _RAND_2952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2953 = {1{`RANDOM}};
  _T_1656_re = _RAND_2953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2954 = {1{`RANDOM}};
  _T_1656_im = _RAND_2954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2955 = {1{`RANDOM}};
  _T_1657_re = _RAND_2955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2956 = {1{`RANDOM}};
  _T_1657_im = _RAND_2956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2957 = {1{`RANDOM}};
  _T_1658_re = _RAND_2957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2958 = {1{`RANDOM}};
  _T_1658_im = _RAND_2958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2959 = {1{`RANDOM}};
  _T_1659_re = _RAND_2959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2960 = {1{`RANDOM}};
  _T_1659_im = _RAND_2960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2961 = {1{`RANDOM}};
  _T_1660_re = _RAND_2961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2962 = {1{`RANDOM}};
  _T_1660_im = _RAND_2962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2963 = {1{`RANDOM}};
  _T_1661_re = _RAND_2963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2964 = {1{`RANDOM}};
  _T_1661_im = _RAND_2964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2965 = {1{`RANDOM}};
  _T_1662_re = _RAND_2965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2966 = {1{`RANDOM}};
  _T_1662_im = _RAND_2966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2967 = {1{`RANDOM}};
  _T_1663_re = _RAND_2967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2968 = {1{`RANDOM}};
  _T_1663_im = _RAND_2968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2969 = {1{`RANDOM}};
  _T_1664_re = _RAND_2969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2970 = {1{`RANDOM}};
  _T_1664_im = _RAND_2970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2971 = {1{`RANDOM}};
  _T_1665_re = _RAND_2971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2972 = {1{`RANDOM}};
  _T_1665_im = _RAND_2972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2973 = {1{`RANDOM}};
  _T_1666_re = _RAND_2973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2974 = {1{`RANDOM}};
  _T_1666_im = _RAND_2974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2975 = {1{`RANDOM}};
  _T_1667_re = _RAND_2975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2976 = {1{`RANDOM}};
  _T_1667_im = _RAND_2976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2977 = {1{`RANDOM}};
  _T_1668_re = _RAND_2977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2978 = {1{`RANDOM}};
  _T_1668_im = _RAND_2978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2979 = {1{`RANDOM}};
  _T_1669_re = _RAND_2979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2980 = {1{`RANDOM}};
  _T_1669_im = _RAND_2980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2981 = {1{`RANDOM}};
  _T_1670_re = _RAND_2981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2982 = {1{`RANDOM}};
  _T_1670_im = _RAND_2982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2983 = {1{`RANDOM}};
  _T_1671_re = _RAND_2983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2984 = {1{`RANDOM}};
  _T_1671_im = _RAND_2984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2985 = {1{`RANDOM}};
  _T_1672_re = _RAND_2985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2986 = {1{`RANDOM}};
  _T_1672_im = _RAND_2986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2987 = {1{`RANDOM}};
  _T_1673_re = _RAND_2987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2988 = {1{`RANDOM}};
  _T_1673_im = _RAND_2988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2989 = {1{`RANDOM}};
  _T_1674_re = _RAND_2989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2990 = {1{`RANDOM}};
  _T_1674_im = _RAND_2990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2991 = {1{`RANDOM}};
  _T_1675_re = _RAND_2991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2992 = {1{`RANDOM}};
  _T_1675_im = _RAND_2992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2993 = {1{`RANDOM}};
  _T_1676_re = _RAND_2993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2994 = {1{`RANDOM}};
  _T_1676_im = _RAND_2994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2995 = {1{`RANDOM}};
  _T_1677_re = _RAND_2995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2996 = {1{`RANDOM}};
  _T_1677_im = _RAND_2996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2997 = {1{`RANDOM}};
  _T_1678_re = _RAND_2997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2998 = {1{`RANDOM}};
  _T_1678_im = _RAND_2998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2999 = {1{`RANDOM}};
  _T_1679_re = _RAND_2999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3000 = {1{`RANDOM}};
  _T_1679_im = _RAND_3000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3001 = {1{`RANDOM}};
  _T_1680_re = _RAND_3001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3002 = {1{`RANDOM}};
  _T_1680_im = _RAND_3002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3003 = {1{`RANDOM}};
  _T_1681_re = _RAND_3003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3004 = {1{`RANDOM}};
  _T_1681_im = _RAND_3004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3005 = {1{`RANDOM}};
  _T_1682_re = _RAND_3005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3006 = {1{`RANDOM}};
  _T_1682_im = _RAND_3006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3007 = {1{`RANDOM}};
  _T_1683_re = _RAND_3007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3008 = {1{`RANDOM}};
  _T_1683_im = _RAND_3008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3009 = {1{`RANDOM}};
  _T_1684_re = _RAND_3009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3010 = {1{`RANDOM}};
  _T_1684_im = _RAND_3010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3011 = {1{`RANDOM}};
  _T_1685_re = _RAND_3011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3012 = {1{`RANDOM}};
  _T_1685_im = _RAND_3012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3013 = {1{`RANDOM}};
  _T_1686_re = _RAND_3013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3014 = {1{`RANDOM}};
  _T_1686_im = _RAND_3014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3015 = {1{`RANDOM}};
  _T_1687_re = _RAND_3015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3016 = {1{`RANDOM}};
  _T_1687_im = _RAND_3016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3017 = {1{`RANDOM}};
  _T_1688_re = _RAND_3017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3018 = {1{`RANDOM}};
  _T_1688_im = _RAND_3018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3019 = {1{`RANDOM}};
  _T_1689_re = _RAND_3019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3020 = {1{`RANDOM}};
  _T_1689_im = _RAND_3020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3021 = {1{`RANDOM}};
  _T_1690_re = _RAND_3021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3022 = {1{`RANDOM}};
  _T_1690_im = _RAND_3022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3023 = {1{`RANDOM}};
  _T_1691_re = _RAND_3023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3024 = {1{`RANDOM}};
  _T_1691_im = _RAND_3024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3025 = {1{`RANDOM}};
  _T_1692_re = _RAND_3025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3026 = {1{`RANDOM}};
  _T_1692_im = _RAND_3026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3027 = {1{`RANDOM}};
  _T_1693_re = _RAND_3027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3028 = {1{`RANDOM}};
  _T_1693_im = _RAND_3028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3029 = {1{`RANDOM}};
  _T_1694_re = _RAND_3029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3030 = {1{`RANDOM}};
  _T_1694_im = _RAND_3030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3031 = {1{`RANDOM}};
  _T_1695_re = _RAND_3031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3032 = {1{`RANDOM}};
  _T_1695_im = _RAND_3032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3033 = {1{`RANDOM}};
  _T_1696_re = _RAND_3033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3034 = {1{`RANDOM}};
  _T_1696_im = _RAND_3034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3035 = {1{`RANDOM}};
  _T_1697_re = _RAND_3035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3036 = {1{`RANDOM}};
  _T_1697_im = _RAND_3036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3037 = {1{`RANDOM}};
  _T_1698_re = _RAND_3037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3038 = {1{`RANDOM}};
  _T_1698_im = _RAND_3038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3039 = {1{`RANDOM}};
  _T_1699_re = _RAND_3039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3040 = {1{`RANDOM}};
  _T_1699_im = _RAND_3040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3041 = {1{`RANDOM}};
  _T_1700_re = _RAND_3041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3042 = {1{`RANDOM}};
  _T_1700_im = _RAND_3042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3043 = {1{`RANDOM}};
  _T_1701_re = _RAND_3043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3044 = {1{`RANDOM}};
  _T_1701_im = _RAND_3044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3045 = {1{`RANDOM}};
  _T_1702_re = _RAND_3045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3046 = {1{`RANDOM}};
  _T_1702_im = _RAND_3046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3047 = {1{`RANDOM}};
  _T_1703_re = _RAND_3047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3048 = {1{`RANDOM}};
  _T_1703_im = _RAND_3048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3049 = {1{`RANDOM}};
  _T_1704_re = _RAND_3049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3050 = {1{`RANDOM}};
  _T_1704_im = _RAND_3050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3051 = {1{`RANDOM}};
  _T_1705_re = _RAND_3051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3052 = {1{`RANDOM}};
  _T_1705_im = _RAND_3052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3053 = {1{`RANDOM}};
  _T_1706_re = _RAND_3053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3054 = {1{`RANDOM}};
  _T_1706_im = _RAND_3054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3055 = {1{`RANDOM}};
  _T_1707_re = _RAND_3055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3056 = {1{`RANDOM}};
  _T_1707_im = _RAND_3056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3057 = {1{`RANDOM}};
  _T_1708_re = _RAND_3057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3058 = {1{`RANDOM}};
  _T_1708_im = _RAND_3058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3059 = {1{`RANDOM}};
  _T_1709_re = _RAND_3059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3060 = {1{`RANDOM}};
  _T_1709_im = _RAND_3060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3061 = {1{`RANDOM}};
  _T_1710_re = _RAND_3061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3062 = {1{`RANDOM}};
  _T_1710_im = _RAND_3062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3063 = {1{`RANDOM}};
  _T_1711_re = _RAND_3063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3064 = {1{`RANDOM}};
  _T_1711_im = _RAND_3064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3065 = {1{`RANDOM}};
  _T_1712_re = _RAND_3065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3066 = {1{`RANDOM}};
  _T_1712_im = _RAND_3066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3067 = {1{`RANDOM}};
  _T_1713_re = _RAND_3067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3068 = {1{`RANDOM}};
  _T_1713_im = _RAND_3068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3069 = {1{`RANDOM}};
  _T_1714_re = _RAND_3069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3070 = {1{`RANDOM}};
  _T_1714_im = _RAND_3070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3071 = {1{`RANDOM}};
  _T_1715_re = _RAND_3071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3072 = {1{`RANDOM}};
  _T_1715_im = _RAND_3072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3073 = {1{`RANDOM}};
  _T_1716_re = _RAND_3073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3074 = {1{`RANDOM}};
  _T_1716_im = _RAND_3074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3075 = {1{`RANDOM}};
  _T_1717_re = _RAND_3075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3076 = {1{`RANDOM}};
  _T_1717_im = _RAND_3076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3077 = {1{`RANDOM}};
  _T_1718_re = _RAND_3077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3078 = {1{`RANDOM}};
  _T_1718_im = _RAND_3078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3079 = {1{`RANDOM}};
  _T_1728_re = _RAND_3079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3080 = {1{`RANDOM}};
  _T_1728_im = _RAND_3080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3081 = {1{`RANDOM}};
  _T_1729_re = _RAND_3081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3082 = {1{`RANDOM}};
  _T_1729_im = _RAND_3082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3083 = {1{`RANDOM}};
  _T_1730_re = _RAND_3083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3084 = {1{`RANDOM}};
  _T_1730_im = _RAND_3084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3085 = {1{`RANDOM}};
  _T_1731_re = _RAND_3085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3086 = {1{`RANDOM}};
  _T_1731_im = _RAND_3086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3087 = {1{`RANDOM}};
  _T_1732_re = _RAND_3087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3088 = {1{`RANDOM}};
  _T_1732_im = _RAND_3088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3089 = {1{`RANDOM}};
  _T_1733_re = _RAND_3089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3090 = {1{`RANDOM}};
  _T_1733_im = _RAND_3090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3091 = {1{`RANDOM}};
  _T_1734_re = _RAND_3091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3092 = {1{`RANDOM}};
  _T_1734_im = _RAND_3092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3093 = {1{`RANDOM}};
  _T_1735_re = _RAND_3093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3094 = {1{`RANDOM}};
  _T_1735_im = _RAND_3094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3095 = {1{`RANDOM}};
  _T_1736_re = _RAND_3095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3096 = {1{`RANDOM}};
  _T_1736_im = _RAND_3096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3097 = {1{`RANDOM}};
  _T_1737_re = _RAND_3097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3098 = {1{`RANDOM}};
  _T_1737_im = _RAND_3098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3099 = {1{`RANDOM}};
  _T_1738_re = _RAND_3099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3100 = {1{`RANDOM}};
  _T_1738_im = _RAND_3100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3101 = {1{`RANDOM}};
  _T_1739_re = _RAND_3101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3102 = {1{`RANDOM}};
  _T_1739_im = _RAND_3102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3103 = {1{`RANDOM}};
  _T_1740_re = _RAND_3103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3104 = {1{`RANDOM}};
  _T_1740_im = _RAND_3104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3105 = {1{`RANDOM}};
  _T_1741_re = _RAND_3105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3106 = {1{`RANDOM}};
  _T_1741_im = _RAND_3106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3107 = {1{`RANDOM}};
  _T_1742_re = _RAND_3107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3108 = {1{`RANDOM}};
  _T_1742_im = _RAND_3108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3109 = {1{`RANDOM}};
  _T_1743_re = _RAND_3109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3110 = {1{`RANDOM}};
  _T_1743_im = _RAND_3110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3111 = {1{`RANDOM}};
  _T_1744_re = _RAND_3111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3112 = {1{`RANDOM}};
  _T_1744_im = _RAND_3112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3113 = {1{`RANDOM}};
  _T_1745_re = _RAND_3113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3114 = {1{`RANDOM}};
  _T_1745_im = _RAND_3114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3115 = {1{`RANDOM}};
  _T_1746_re = _RAND_3115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3116 = {1{`RANDOM}};
  _T_1746_im = _RAND_3116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3117 = {1{`RANDOM}};
  _T_1747_re = _RAND_3117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3118 = {1{`RANDOM}};
  _T_1747_im = _RAND_3118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3119 = {1{`RANDOM}};
  _T_1748_re = _RAND_3119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3120 = {1{`RANDOM}};
  _T_1748_im = _RAND_3120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3121 = {1{`RANDOM}};
  _T_1749_re = _RAND_3121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3122 = {1{`RANDOM}};
  _T_1749_im = _RAND_3122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3123 = {1{`RANDOM}};
  _T_1750_re = _RAND_3123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3124 = {1{`RANDOM}};
  _T_1750_im = _RAND_3124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3125 = {1{`RANDOM}};
  _T_1751_re = _RAND_3125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3126 = {1{`RANDOM}};
  _T_1751_im = _RAND_3126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3127 = {1{`RANDOM}};
  _T_1752_re = _RAND_3127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3128 = {1{`RANDOM}};
  _T_1752_im = _RAND_3128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3129 = {1{`RANDOM}};
  _T_1753_re = _RAND_3129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3130 = {1{`RANDOM}};
  _T_1753_im = _RAND_3130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3131 = {1{`RANDOM}};
  _T_1754_re = _RAND_3131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3132 = {1{`RANDOM}};
  _T_1754_im = _RAND_3132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3133 = {1{`RANDOM}};
  _T_1755_re = _RAND_3133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3134 = {1{`RANDOM}};
  _T_1755_im = _RAND_3134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3135 = {1{`RANDOM}};
  _T_1756_re = _RAND_3135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3136 = {1{`RANDOM}};
  _T_1756_im = _RAND_3136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3137 = {1{`RANDOM}};
  _T_1757_re = _RAND_3137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3138 = {1{`RANDOM}};
  _T_1757_im = _RAND_3138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3139 = {1{`RANDOM}};
  _T_1758_re = _RAND_3139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3140 = {1{`RANDOM}};
  _T_1758_im = _RAND_3140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3141 = {1{`RANDOM}};
  _T_1759_re = _RAND_3141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3142 = {1{`RANDOM}};
  _T_1759_im = _RAND_3142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3143 = {1{`RANDOM}};
  _T_1760_re = _RAND_3143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3144 = {1{`RANDOM}};
  _T_1760_im = _RAND_3144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3145 = {1{`RANDOM}};
  _T_1761_re = _RAND_3145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3146 = {1{`RANDOM}};
  _T_1761_im = _RAND_3146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3147 = {1{`RANDOM}};
  _T_1762_re = _RAND_3147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3148 = {1{`RANDOM}};
  _T_1762_im = _RAND_3148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3149 = {1{`RANDOM}};
  _T_1763_re = _RAND_3149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3150 = {1{`RANDOM}};
  _T_1763_im = _RAND_3150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3151 = {1{`RANDOM}};
  _T_1764_re = _RAND_3151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3152 = {1{`RANDOM}};
  _T_1764_im = _RAND_3152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3153 = {1{`RANDOM}};
  _T_1765_re = _RAND_3153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3154 = {1{`RANDOM}};
  _T_1765_im = _RAND_3154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3155 = {1{`RANDOM}};
  _T_1766_re = _RAND_3155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3156 = {1{`RANDOM}};
  _T_1766_im = _RAND_3156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3157 = {1{`RANDOM}};
  _T_1767_re = _RAND_3157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3158 = {1{`RANDOM}};
  _T_1767_im = _RAND_3158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3159 = {1{`RANDOM}};
  _T_1768_re = _RAND_3159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3160 = {1{`RANDOM}};
  _T_1768_im = _RAND_3160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3161 = {1{`RANDOM}};
  _T_1769_re = _RAND_3161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3162 = {1{`RANDOM}};
  _T_1769_im = _RAND_3162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3163 = {1{`RANDOM}};
  _T_1770_re = _RAND_3163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3164 = {1{`RANDOM}};
  _T_1770_im = _RAND_3164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3165 = {1{`RANDOM}};
  _T_1771_re = _RAND_3165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3166 = {1{`RANDOM}};
  _T_1771_im = _RAND_3166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3167 = {1{`RANDOM}};
  _T_1772_re = _RAND_3167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3168 = {1{`RANDOM}};
  _T_1772_im = _RAND_3168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3169 = {1{`RANDOM}};
  _T_1773_re = _RAND_3169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3170 = {1{`RANDOM}};
  _T_1773_im = _RAND_3170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3171 = {1{`RANDOM}};
  _T_1774_re = _RAND_3171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3172 = {1{`RANDOM}};
  _T_1774_im = _RAND_3172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3173 = {1{`RANDOM}};
  _T_1775_re = _RAND_3173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3174 = {1{`RANDOM}};
  _T_1775_im = _RAND_3174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3175 = {1{`RANDOM}};
  _T_1776_re = _RAND_3175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3176 = {1{`RANDOM}};
  _T_1776_im = _RAND_3176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3177 = {1{`RANDOM}};
  _T_1777_re = _RAND_3177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3178 = {1{`RANDOM}};
  _T_1777_im = _RAND_3178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3179 = {1{`RANDOM}};
  _T_1778_re = _RAND_3179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3180 = {1{`RANDOM}};
  _T_1778_im = _RAND_3180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3181 = {1{`RANDOM}};
  _T_1779_re = _RAND_3181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3182 = {1{`RANDOM}};
  _T_1779_im = _RAND_3182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3183 = {1{`RANDOM}};
  _T_1780_re = _RAND_3183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3184 = {1{`RANDOM}};
  _T_1780_im = _RAND_3184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3185 = {1{`RANDOM}};
  _T_1781_re = _RAND_3185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3186 = {1{`RANDOM}};
  _T_1781_im = _RAND_3186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3187 = {1{`RANDOM}};
  _T_1782_re = _RAND_3187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3188 = {1{`RANDOM}};
  _T_1782_im = _RAND_3188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3189 = {1{`RANDOM}};
  _T_1783_re = _RAND_3189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3190 = {1{`RANDOM}};
  _T_1783_im = _RAND_3190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3191 = {1{`RANDOM}};
  _T_1784_re = _RAND_3191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3192 = {1{`RANDOM}};
  _T_1784_im = _RAND_3192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3193 = {1{`RANDOM}};
  _T_1785_re = _RAND_3193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3194 = {1{`RANDOM}};
  _T_1785_im = _RAND_3194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3195 = {1{`RANDOM}};
  _T_1786_re = _RAND_3195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3196 = {1{`RANDOM}};
  _T_1786_im = _RAND_3196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3197 = {1{`RANDOM}};
  _T_1787_re = _RAND_3197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3198 = {1{`RANDOM}};
  _T_1787_im = _RAND_3198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3199 = {1{`RANDOM}};
  _T_1788_re = _RAND_3199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3200 = {1{`RANDOM}};
  _T_1788_im = _RAND_3200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3201 = {1{`RANDOM}};
  _T_1789_re = _RAND_3201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3202 = {1{`RANDOM}};
  _T_1789_im = _RAND_3202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3203 = {1{`RANDOM}};
  _T_1790_re = _RAND_3203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3204 = {1{`RANDOM}};
  _T_1790_im = _RAND_3204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3205 = {1{`RANDOM}};
  _T_1791_re = _RAND_3205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3206 = {1{`RANDOM}};
  _T_1791_im = _RAND_3206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3207 = {1{`RANDOM}};
  _T_1792_re = _RAND_3207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3208 = {1{`RANDOM}};
  _T_1792_im = _RAND_3208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3209 = {1{`RANDOM}};
  _T_1793_re = _RAND_3209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3210 = {1{`RANDOM}};
  _T_1793_im = _RAND_3210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3211 = {1{`RANDOM}};
  _T_1794_re = _RAND_3211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3212 = {1{`RANDOM}};
  _T_1794_im = _RAND_3212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3213 = {1{`RANDOM}};
  _T_1795_re = _RAND_3213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3214 = {1{`RANDOM}};
  _T_1795_im = _RAND_3214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3215 = {1{`RANDOM}};
  _T_1796_re = _RAND_3215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3216 = {1{`RANDOM}};
  _T_1796_im = _RAND_3216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3217 = {1{`RANDOM}};
  _T_1797_re = _RAND_3217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3218 = {1{`RANDOM}};
  _T_1797_im = _RAND_3218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3219 = {1{`RANDOM}};
  _T_1798_re = _RAND_3219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3220 = {1{`RANDOM}};
  _T_1798_im = _RAND_3220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3221 = {1{`RANDOM}};
  _T_1799_re = _RAND_3221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3222 = {1{`RANDOM}};
  _T_1799_im = _RAND_3222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3223 = {1{`RANDOM}};
  _T_1800_re = _RAND_3223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3224 = {1{`RANDOM}};
  _T_1800_im = _RAND_3224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3225 = {1{`RANDOM}};
  _T_1801_re = _RAND_3225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3226 = {1{`RANDOM}};
  _T_1801_im = _RAND_3226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3227 = {1{`RANDOM}};
  _T_1802_re = _RAND_3227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3228 = {1{`RANDOM}};
  _T_1802_im = _RAND_3228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3229 = {1{`RANDOM}};
  _T_1803_re = _RAND_3229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3230 = {1{`RANDOM}};
  _T_1803_im = _RAND_3230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3231 = {1{`RANDOM}};
  _T_1804_re = _RAND_3231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3232 = {1{`RANDOM}};
  _T_1804_im = _RAND_3232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3233 = {1{`RANDOM}};
  _T_1805_re = _RAND_3233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3234 = {1{`RANDOM}};
  _T_1805_im = _RAND_3234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3235 = {1{`RANDOM}};
  _T_1806_re = _RAND_3235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3236 = {1{`RANDOM}};
  _T_1806_im = _RAND_3236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3237 = {1{`RANDOM}};
  _T_1807_re = _RAND_3237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3238 = {1{`RANDOM}};
  _T_1807_im = _RAND_3238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3239 = {1{`RANDOM}};
  _T_1808_re = _RAND_3239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3240 = {1{`RANDOM}};
  _T_1808_im = _RAND_3240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3241 = {1{`RANDOM}};
  _T_1809_re = _RAND_3241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3242 = {1{`RANDOM}};
  _T_1809_im = _RAND_3242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3243 = {1{`RANDOM}};
  _T_1810_re = _RAND_3243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3244 = {1{`RANDOM}};
  _T_1810_im = _RAND_3244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3245 = {1{`RANDOM}};
  _T_1811_re = _RAND_3245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3246 = {1{`RANDOM}};
  _T_1811_im = _RAND_3246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3247 = {1{`RANDOM}};
  _T_1812_re = _RAND_3247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3248 = {1{`RANDOM}};
  _T_1812_im = _RAND_3248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3249 = {1{`RANDOM}};
  _T_1813_re = _RAND_3249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3250 = {1{`RANDOM}};
  _T_1813_im = _RAND_3250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3251 = {1{`RANDOM}};
  _T_1814_re = _RAND_3251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3252 = {1{`RANDOM}};
  _T_1814_im = _RAND_3252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3253 = {1{`RANDOM}};
  _T_1815_re = _RAND_3253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3254 = {1{`RANDOM}};
  _T_1815_im = _RAND_3254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3255 = {1{`RANDOM}};
  _T_1816_re = _RAND_3255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3256 = {1{`RANDOM}};
  _T_1816_im = _RAND_3256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3257 = {1{`RANDOM}};
  _T_1817_re = _RAND_3257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3258 = {1{`RANDOM}};
  _T_1817_im = _RAND_3258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3259 = {1{`RANDOM}};
  _T_1818_re = _RAND_3259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3260 = {1{`RANDOM}};
  _T_1818_im = _RAND_3260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3261 = {1{`RANDOM}};
  _T_1819_re = _RAND_3261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3262 = {1{`RANDOM}};
  _T_1819_im = _RAND_3262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3263 = {1{`RANDOM}};
  _T_1820_re = _RAND_3263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3264 = {1{`RANDOM}};
  _T_1820_im = _RAND_3264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3265 = {1{`RANDOM}};
  _T_1821_re = _RAND_3265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3266 = {1{`RANDOM}};
  _T_1821_im = _RAND_3266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3267 = {1{`RANDOM}};
  _T_1822_re = _RAND_3267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3268 = {1{`RANDOM}};
  _T_1822_im = _RAND_3268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3269 = {1{`RANDOM}};
  _T_1823_re = _RAND_3269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3270 = {1{`RANDOM}};
  _T_1823_im = _RAND_3270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3271 = {1{`RANDOM}};
  _T_1824_re = _RAND_3271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3272 = {1{`RANDOM}};
  _T_1824_im = _RAND_3272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3273 = {1{`RANDOM}};
  _T_1825_re = _RAND_3273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3274 = {1{`RANDOM}};
  _T_1825_im = _RAND_3274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3275 = {1{`RANDOM}};
  _T_1826_re = _RAND_3275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3276 = {1{`RANDOM}};
  _T_1826_im = _RAND_3276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3277 = {1{`RANDOM}};
  _T_1827_re = _RAND_3277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3278 = {1{`RANDOM}};
  _T_1827_im = _RAND_3278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3279 = {1{`RANDOM}};
  _T_1828_re = _RAND_3279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3280 = {1{`RANDOM}};
  _T_1828_im = _RAND_3280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3281 = {1{`RANDOM}};
  _T_1829_re = _RAND_3281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3282 = {1{`RANDOM}};
  _T_1829_im = _RAND_3282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3283 = {1{`RANDOM}};
  _T_1830_re = _RAND_3283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3284 = {1{`RANDOM}};
  _T_1830_im = _RAND_3284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3285 = {1{`RANDOM}};
  _T_1831_re = _RAND_3285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3286 = {1{`RANDOM}};
  _T_1831_im = _RAND_3286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3287 = {1{`RANDOM}};
  _T_1832_re = _RAND_3287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3288 = {1{`RANDOM}};
  _T_1832_im = _RAND_3288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3289 = {1{`RANDOM}};
  _T_1833_re = _RAND_3289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3290 = {1{`RANDOM}};
  _T_1833_im = _RAND_3290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3291 = {1{`RANDOM}};
  _T_1834_re = _RAND_3291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3292 = {1{`RANDOM}};
  _T_1834_im = _RAND_3292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3293 = {1{`RANDOM}};
  _T_1835_re = _RAND_3293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3294 = {1{`RANDOM}};
  _T_1835_im = _RAND_3294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3295 = {1{`RANDOM}};
  _T_1836_re = _RAND_3295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3296 = {1{`RANDOM}};
  _T_1836_im = _RAND_3296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3297 = {1{`RANDOM}};
  _T_1837_re = _RAND_3297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3298 = {1{`RANDOM}};
  _T_1837_im = _RAND_3298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3299 = {1{`RANDOM}};
  _T_1838_re = _RAND_3299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3300 = {1{`RANDOM}};
  _T_1838_im = _RAND_3300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3301 = {1{`RANDOM}};
  _T_1839_re = _RAND_3301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3302 = {1{`RANDOM}};
  _T_1839_im = _RAND_3302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3303 = {1{`RANDOM}};
  _T_1840_re = _RAND_3303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3304 = {1{`RANDOM}};
  _T_1840_im = _RAND_3304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3305 = {1{`RANDOM}};
  _T_1841_re = _RAND_3305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3306 = {1{`RANDOM}};
  _T_1841_im = _RAND_3306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3307 = {1{`RANDOM}};
  _T_1842_re = _RAND_3307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3308 = {1{`RANDOM}};
  _T_1842_im = _RAND_3308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3309 = {1{`RANDOM}};
  _T_1843_re = _RAND_3309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3310 = {1{`RANDOM}};
  _T_1843_im = _RAND_3310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3311 = {1{`RANDOM}};
  _T_1844_re = _RAND_3311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3312 = {1{`RANDOM}};
  _T_1844_im = _RAND_3312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3313 = {1{`RANDOM}};
  _T_1845_re = _RAND_3313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3314 = {1{`RANDOM}};
  _T_1845_im = _RAND_3314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3315 = {1{`RANDOM}};
  _T_1846_re = _RAND_3315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3316 = {1{`RANDOM}};
  _T_1846_im = _RAND_3316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3317 = {1{`RANDOM}};
  _T_1847_re = _RAND_3317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3318 = {1{`RANDOM}};
  _T_1847_im = _RAND_3318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3319 = {1{`RANDOM}};
  _T_1848_re = _RAND_3319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3320 = {1{`RANDOM}};
  _T_1848_im = _RAND_3320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3321 = {1{`RANDOM}};
  _T_1849_re = _RAND_3321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3322 = {1{`RANDOM}};
  _T_1849_im = _RAND_3322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3323 = {1{`RANDOM}};
  _T_1850_re = _RAND_3323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3324 = {1{`RANDOM}};
  _T_1850_im = _RAND_3324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3325 = {1{`RANDOM}};
  _T_1851_re = _RAND_3325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3326 = {1{`RANDOM}};
  _T_1851_im = _RAND_3326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3327 = {1{`RANDOM}};
  _T_1852_re = _RAND_3327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3328 = {1{`RANDOM}};
  _T_1852_im = _RAND_3328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3329 = {1{`RANDOM}};
  _T_1853_re = _RAND_3329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3330 = {1{`RANDOM}};
  _T_1853_im = _RAND_3330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3331 = {1{`RANDOM}};
  _T_1854_re = _RAND_3331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3332 = {1{`RANDOM}};
  _T_1854_im = _RAND_3332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3333 = {1{`RANDOM}};
  _T_1855_re = _RAND_3333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3334 = {1{`RANDOM}};
  _T_1855_im = _RAND_3334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3335 = {1{`RANDOM}};
  _T_1856_re = _RAND_3335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3336 = {1{`RANDOM}};
  _T_1856_im = _RAND_3336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3337 = {1{`RANDOM}};
  _T_1857_re = _RAND_3337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3338 = {1{`RANDOM}};
  _T_1857_im = _RAND_3338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3339 = {1{`RANDOM}};
  _T_1858_re = _RAND_3339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3340 = {1{`RANDOM}};
  _T_1858_im = _RAND_3340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3341 = {1{`RANDOM}};
  _T_1859_re = _RAND_3341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3342 = {1{`RANDOM}};
  _T_1859_im = _RAND_3342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3343 = {1{`RANDOM}};
  _T_1860_re = _RAND_3343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3344 = {1{`RANDOM}};
  _T_1860_im = _RAND_3344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3345 = {1{`RANDOM}};
  _T_1861_re = _RAND_3345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3346 = {1{`RANDOM}};
  _T_1861_im = _RAND_3346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3347 = {1{`RANDOM}};
  _T_1862_re = _RAND_3347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3348 = {1{`RANDOM}};
  _T_1862_im = _RAND_3348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3349 = {1{`RANDOM}};
  _T_1863_re = _RAND_3349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3350 = {1{`RANDOM}};
  _T_1863_im = _RAND_3350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3351 = {1{`RANDOM}};
  _T_1864_re = _RAND_3351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3352 = {1{`RANDOM}};
  _T_1864_im = _RAND_3352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3353 = {1{`RANDOM}};
  _T_1865_re = _RAND_3353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3354 = {1{`RANDOM}};
  _T_1865_im = _RAND_3354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3355 = {1{`RANDOM}};
  _T_1866_re = _RAND_3355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3356 = {1{`RANDOM}};
  _T_1866_im = _RAND_3356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3357 = {1{`RANDOM}};
  _T_1867_re = _RAND_3357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3358 = {1{`RANDOM}};
  _T_1867_im = _RAND_3358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3359 = {1{`RANDOM}};
  _T_1868_re = _RAND_3359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3360 = {1{`RANDOM}};
  _T_1868_im = _RAND_3360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3361 = {1{`RANDOM}};
  _T_1869_re = _RAND_3361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3362 = {1{`RANDOM}};
  _T_1869_im = _RAND_3362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3363 = {1{`RANDOM}};
  _T_1870_re = _RAND_3363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3364 = {1{`RANDOM}};
  _T_1870_im = _RAND_3364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3365 = {1{`RANDOM}};
  _T_1871_re = _RAND_3365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3366 = {1{`RANDOM}};
  _T_1871_im = _RAND_3366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3367 = {1{`RANDOM}};
  _T_1872_re = _RAND_3367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3368 = {1{`RANDOM}};
  _T_1872_im = _RAND_3368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3369 = {1{`RANDOM}};
  _T_1873_re = _RAND_3369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3370 = {1{`RANDOM}};
  _T_1873_im = _RAND_3370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3371 = {1{`RANDOM}};
  _T_1874_re = _RAND_3371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3372 = {1{`RANDOM}};
  _T_1874_im = _RAND_3372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3373 = {1{`RANDOM}};
  _T_1875_re = _RAND_3373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3374 = {1{`RANDOM}};
  _T_1875_im = _RAND_3374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3375 = {1{`RANDOM}};
  _T_1876_re = _RAND_3375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3376 = {1{`RANDOM}};
  _T_1876_im = _RAND_3376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3377 = {1{`RANDOM}};
  _T_1877_re = _RAND_3377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3378 = {1{`RANDOM}};
  _T_1877_im = _RAND_3378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3379 = {1{`RANDOM}};
  _T_1878_re = _RAND_3379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3380 = {1{`RANDOM}};
  _T_1878_im = _RAND_3380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3381 = {1{`RANDOM}};
  _T_1879_re = _RAND_3381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3382 = {1{`RANDOM}};
  _T_1879_im = _RAND_3382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3383 = {1{`RANDOM}};
  _T_1880_re = _RAND_3383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3384 = {1{`RANDOM}};
  _T_1880_im = _RAND_3384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3385 = {1{`RANDOM}};
  _T_1881_re = _RAND_3385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3386 = {1{`RANDOM}};
  _T_1881_im = _RAND_3386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3387 = {1{`RANDOM}};
  _T_1882_re = _RAND_3387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3388 = {1{`RANDOM}};
  _T_1882_im = _RAND_3388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3389 = {1{`RANDOM}};
  _T_1883_re = _RAND_3389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3390 = {1{`RANDOM}};
  _T_1883_im = _RAND_3390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3391 = {1{`RANDOM}};
  _T_1884_re = _RAND_3391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3392 = {1{`RANDOM}};
  _T_1884_im = _RAND_3392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3393 = {1{`RANDOM}};
  _T_1885_re = _RAND_3393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3394 = {1{`RANDOM}};
  _T_1885_im = _RAND_3394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3395 = {1{`RANDOM}};
  _T_1886_re = _RAND_3395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3396 = {1{`RANDOM}};
  _T_1886_im = _RAND_3396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3397 = {1{`RANDOM}};
  _T_1887_re = _RAND_3397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3398 = {1{`RANDOM}};
  _T_1887_im = _RAND_3398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3399 = {1{`RANDOM}};
  _T_1888_re = _RAND_3399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3400 = {1{`RANDOM}};
  _T_1888_im = _RAND_3400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3401 = {1{`RANDOM}};
  _T_1889_re = _RAND_3401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3402 = {1{`RANDOM}};
  _T_1889_im = _RAND_3402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3403 = {1{`RANDOM}};
  _T_1890_re = _RAND_3403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3404 = {1{`RANDOM}};
  _T_1890_im = _RAND_3404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3405 = {1{`RANDOM}};
  _T_1891_re = _RAND_3405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3406 = {1{`RANDOM}};
  _T_1891_im = _RAND_3406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3407 = {1{`RANDOM}};
  _T_1892_re = _RAND_3407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3408 = {1{`RANDOM}};
  _T_1892_im = _RAND_3408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3409 = {1{`RANDOM}};
  _T_1893_re = _RAND_3409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3410 = {1{`RANDOM}};
  _T_1893_im = _RAND_3410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3411 = {1{`RANDOM}};
  _T_1894_re = _RAND_3411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3412 = {1{`RANDOM}};
  _T_1894_im = _RAND_3412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3413 = {1{`RANDOM}};
  _T_1895_re = _RAND_3413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3414 = {1{`RANDOM}};
  _T_1895_im = _RAND_3414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3415 = {1{`RANDOM}};
  _T_1896_re = _RAND_3415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3416 = {1{`RANDOM}};
  _T_1896_im = _RAND_3416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3417 = {1{`RANDOM}};
  _T_1897_re = _RAND_3417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3418 = {1{`RANDOM}};
  _T_1897_im = _RAND_3418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3419 = {1{`RANDOM}};
  _T_1898_re = _RAND_3419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3420 = {1{`RANDOM}};
  _T_1898_im = _RAND_3420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3421 = {1{`RANDOM}};
  _T_1899_re = _RAND_3421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3422 = {1{`RANDOM}};
  _T_1899_im = _RAND_3422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3423 = {1{`RANDOM}};
  _T_1900_re = _RAND_3423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3424 = {1{`RANDOM}};
  _T_1900_im = _RAND_3424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3425 = {1{`RANDOM}};
  _T_1901_re = _RAND_3425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3426 = {1{`RANDOM}};
  _T_1901_im = _RAND_3426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3427 = {1{`RANDOM}};
  _T_1902_re = _RAND_3427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3428 = {1{`RANDOM}};
  _T_1902_im = _RAND_3428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3429 = {1{`RANDOM}};
  _T_1903_re = _RAND_3429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3430 = {1{`RANDOM}};
  _T_1903_im = _RAND_3430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3431 = {1{`RANDOM}};
  _T_1904_re = _RAND_3431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3432 = {1{`RANDOM}};
  _T_1904_im = _RAND_3432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3433 = {1{`RANDOM}};
  _T_1905_re = _RAND_3433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3434 = {1{`RANDOM}};
  _T_1905_im = _RAND_3434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3435 = {1{`RANDOM}};
  _T_1906_re = _RAND_3435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3436 = {1{`RANDOM}};
  _T_1906_im = _RAND_3436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3437 = {1{`RANDOM}};
  _T_1907_re = _RAND_3437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3438 = {1{`RANDOM}};
  _T_1907_im = _RAND_3438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3439 = {1{`RANDOM}};
  _T_1908_re = _RAND_3439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3440 = {1{`RANDOM}};
  _T_1908_im = _RAND_3440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3441 = {1{`RANDOM}};
  _T_1909_re = _RAND_3441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3442 = {1{`RANDOM}};
  _T_1909_im = _RAND_3442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3443 = {1{`RANDOM}};
  _T_1910_re = _RAND_3443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3444 = {1{`RANDOM}};
  _T_1910_im = _RAND_3444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3445 = {1{`RANDOM}};
  _T_1911_re = _RAND_3445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3446 = {1{`RANDOM}};
  _T_1911_im = _RAND_3446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3447 = {1{`RANDOM}};
  _T_1912_re = _RAND_3447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3448 = {1{`RANDOM}};
  _T_1912_im = _RAND_3448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3449 = {1{`RANDOM}};
  _T_1913_re = _RAND_3449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3450 = {1{`RANDOM}};
  _T_1913_im = _RAND_3450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3451 = {1{`RANDOM}};
  _T_1914_re = _RAND_3451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3452 = {1{`RANDOM}};
  _T_1914_im = _RAND_3452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3453 = {1{`RANDOM}};
  _T_1915_re = _RAND_3453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3454 = {1{`RANDOM}};
  _T_1915_im = _RAND_3454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3455 = {1{`RANDOM}};
  _T_1916_re = _RAND_3455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3456 = {1{`RANDOM}};
  _T_1916_im = _RAND_3456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3457 = {1{`RANDOM}};
  _T_1917_re = _RAND_3457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3458 = {1{`RANDOM}};
  _T_1917_im = _RAND_3458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3459 = {1{`RANDOM}};
  _T_1918_re = _RAND_3459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3460 = {1{`RANDOM}};
  _T_1918_im = _RAND_3460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3461 = {1{`RANDOM}};
  _T_1919_re = _RAND_3461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3462 = {1{`RANDOM}};
  _T_1919_im = _RAND_3462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3463 = {1{`RANDOM}};
  _T_1920_re = _RAND_3463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3464 = {1{`RANDOM}};
  _T_1920_im = _RAND_3464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3465 = {1{`RANDOM}};
  _T_1921_re = _RAND_3465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3466 = {1{`RANDOM}};
  _T_1921_im = _RAND_3466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3467 = {1{`RANDOM}};
  _T_1922_re = _RAND_3467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3468 = {1{`RANDOM}};
  _T_1922_im = _RAND_3468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3469 = {1{`RANDOM}};
  _T_1923_re = _RAND_3469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3470 = {1{`RANDOM}};
  _T_1923_im = _RAND_3470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3471 = {1{`RANDOM}};
  _T_1924_re = _RAND_3471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3472 = {1{`RANDOM}};
  _T_1924_im = _RAND_3472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3473 = {1{`RANDOM}};
  _T_1925_re = _RAND_3473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3474 = {1{`RANDOM}};
  _T_1925_im = _RAND_3474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3475 = {1{`RANDOM}};
  _T_1926_re = _RAND_3475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3476 = {1{`RANDOM}};
  _T_1926_im = _RAND_3476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3477 = {1{`RANDOM}};
  _T_1927_re = _RAND_3477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3478 = {1{`RANDOM}};
  _T_1927_im = _RAND_3478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3479 = {1{`RANDOM}};
  _T_1928_re = _RAND_3479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3480 = {1{`RANDOM}};
  _T_1928_im = _RAND_3480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3481 = {1{`RANDOM}};
  _T_1929_re = _RAND_3481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3482 = {1{`RANDOM}};
  _T_1929_im = _RAND_3482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3483 = {1{`RANDOM}};
  _T_1930_re = _RAND_3483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3484 = {1{`RANDOM}};
  _T_1930_im = _RAND_3484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3485 = {1{`RANDOM}};
  _T_1931_re = _RAND_3485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3486 = {1{`RANDOM}};
  _T_1931_im = _RAND_3486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3487 = {1{`RANDOM}};
  _T_1932_re = _RAND_3487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3488 = {1{`RANDOM}};
  _T_1932_im = _RAND_3488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3489 = {1{`RANDOM}};
  _T_1933_re = _RAND_3489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3490 = {1{`RANDOM}};
  _T_1933_im = _RAND_3490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3491 = {1{`RANDOM}};
  _T_1934_re = _RAND_3491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3492 = {1{`RANDOM}};
  _T_1934_im = _RAND_3492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3493 = {1{`RANDOM}};
  _T_1935_re = _RAND_3493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3494 = {1{`RANDOM}};
  _T_1935_im = _RAND_3494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3495 = {1{`RANDOM}};
  _T_1936_re = _RAND_3495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3496 = {1{`RANDOM}};
  _T_1936_im = _RAND_3496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3497 = {1{`RANDOM}};
  _T_1937_re = _RAND_3497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3498 = {1{`RANDOM}};
  _T_1937_im = _RAND_3498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3499 = {1{`RANDOM}};
  _T_1938_re = _RAND_3499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3500 = {1{`RANDOM}};
  _T_1938_im = _RAND_3500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3501 = {1{`RANDOM}};
  _T_1939_re = _RAND_3501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3502 = {1{`RANDOM}};
  _T_1939_im = _RAND_3502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3503 = {1{`RANDOM}};
  _T_1940_re = _RAND_3503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3504 = {1{`RANDOM}};
  _T_1940_im = _RAND_3504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3505 = {1{`RANDOM}};
  _T_1941_re = _RAND_3505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3506 = {1{`RANDOM}};
  _T_1941_im = _RAND_3506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3507 = {1{`RANDOM}};
  _T_1942_re = _RAND_3507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3508 = {1{`RANDOM}};
  _T_1942_im = _RAND_3508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3509 = {1{`RANDOM}};
  _T_1943_re = _RAND_3509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3510 = {1{`RANDOM}};
  _T_1943_im = _RAND_3510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3511 = {1{`RANDOM}};
  _T_1944_re = _RAND_3511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3512 = {1{`RANDOM}};
  _T_1944_im = _RAND_3512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3513 = {1{`RANDOM}};
  _T_1945_re = _RAND_3513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3514 = {1{`RANDOM}};
  _T_1945_im = _RAND_3514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3515 = {1{`RANDOM}};
  _T_1946_re = _RAND_3515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3516 = {1{`RANDOM}};
  _T_1946_im = _RAND_3516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3517 = {1{`RANDOM}};
  _T_1947_re = _RAND_3517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3518 = {1{`RANDOM}};
  _T_1947_im = _RAND_3518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3519 = {1{`RANDOM}};
  _T_1948_re = _RAND_3519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3520 = {1{`RANDOM}};
  _T_1948_im = _RAND_3520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3521 = {1{`RANDOM}};
  _T_1949_re = _RAND_3521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3522 = {1{`RANDOM}};
  _T_1949_im = _RAND_3522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3523 = {1{`RANDOM}};
  _T_1950_re = _RAND_3523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3524 = {1{`RANDOM}};
  _T_1950_im = _RAND_3524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3525 = {1{`RANDOM}};
  _T_1951_re = _RAND_3525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3526 = {1{`RANDOM}};
  _T_1951_im = _RAND_3526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3527 = {1{`RANDOM}};
  _T_1952_re = _RAND_3527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3528 = {1{`RANDOM}};
  _T_1952_im = _RAND_3528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3529 = {1{`RANDOM}};
  _T_1953_re = _RAND_3529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3530 = {1{`RANDOM}};
  _T_1953_im = _RAND_3530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3531 = {1{`RANDOM}};
  _T_1954_re = _RAND_3531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3532 = {1{`RANDOM}};
  _T_1954_im = _RAND_3532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3533 = {1{`RANDOM}};
  _T_1955_re = _RAND_3533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3534 = {1{`RANDOM}};
  _T_1955_im = _RAND_3534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3535 = {1{`RANDOM}};
  _T_1956_re = _RAND_3535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3536 = {1{`RANDOM}};
  _T_1956_im = _RAND_3536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3537 = {1{`RANDOM}};
  _T_1957_re = _RAND_3537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3538 = {1{`RANDOM}};
  _T_1957_im = _RAND_3538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3539 = {1{`RANDOM}};
  _T_1958_re = _RAND_3539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3540 = {1{`RANDOM}};
  _T_1958_im = _RAND_3540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3541 = {1{`RANDOM}};
  _T_1959_re = _RAND_3541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3542 = {1{`RANDOM}};
  _T_1959_im = _RAND_3542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3543 = {1{`RANDOM}};
  _T_1960_re = _RAND_3543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3544 = {1{`RANDOM}};
  _T_1960_im = _RAND_3544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3545 = {1{`RANDOM}};
  _T_1961_re = _RAND_3545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3546 = {1{`RANDOM}};
  _T_1961_im = _RAND_3546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3547 = {1{`RANDOM}};
  _T_1962_re = _RAND_3547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3548 = {1{`RANDOM}};
  _T_1962_im = _RAND_3548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3549 = {1{`RANDOM}};
  _T_1963_re = _RAND_3549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3550 = {1{`RANDOM}};
  _T_1963_im = _RAND_3550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3551 = {1{`RANDOM}};
  _T_1964_re = _RAND_3551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3552 = {1{`RANDOM}};
  _T_1964_im = _RAND_3552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3553 = {1{`RANDOM}};
  _T_1965_re = _RAND_3553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3554 = {1{`RANDOM}};
  _T_1965_im = _RAND_3554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3555 = {1{`RANDOM}};
  _T_1966_re = _RAND_3555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3556 = {1{`RANDOM}};
  _T_1966_im = _RAND_3556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3557 = {1{`RANDOM}};
  _T_1967_re = _RAND_3557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3558 = {1{`RANDOM}};
  _T_1967_im = _RAND_3558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3559 = {1{`RANDOM}};
  _T_1968_re = _RAND_3559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3560 = {1{`RANDOM}};
  _T_1968_im = _RAND_3560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3561 = {1{`RANDOM}};
  _T_1969_re = _RAND_3561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3562 = {1{`RANDOM}};
  _T_1969_im = _RAND_3562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3563 = {1{`RANDOM}};
  _T_1970_re = _RAND_3563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3564 = {1{`RANDOM}};
  _T_1970_im = _RAND_3564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3565 = {1{`RANDOM}};
  _T_1971_re = _RAND_3565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3566 = {1{`RANDOM}};
  _T_1971_im = _RAND_3566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3567 = {1{`RANDOM}};
  _T_1972_re = _RAND_3567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3568 = {1{`RANDOM}};
  _T_1972_im = _RAND_3568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3569 = {1{`RANDOM}};
  _T_1973_re = _RAND_3569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3570 = {1{`RANDOM}};
  _T_1973_im = _RAND_3570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3571 = {1{`RANDOM}};
  _T_1974_re = _RAND_3571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3572 = {1{`RANDOM}};
  _T_1974_im = _RAND_3572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3573 = {1{`RANDOM}};
  _T_1975_re = _RAND_3573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3574 = {1{`RANDOM}};
  _T_1975_im = _RAND_3574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3575 = {1{`RANDOM}};
  _T_1976_re = _RAND_3575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3576 = {1{`RANDOM}};
  _T_1976_im = _RAND_3576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3577 = {1{`RANDOM}};
  _T_1977_re = _RAND_3577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3578 = {1{`RANDOM}};
  _T_1977_im = _RAND_3578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3579 = {1{`RANDOM}};
  _T_1978_re = _RAND_3579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3580 = {1{`RANDOM}};
  _T_1978_im = _RAND_3580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3581 = {1{`RANDOM}};
  _T_1979_re = _RAND_3581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3582 = {1{`RANDOM}};
  _T_1979_im = _RAND_3582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3583 = {1{`RANDOM}};
  _T_1980_re = _RAND_3583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3584 = {1{`RANDOM}};
  _T_1980_im = _RAND_3584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3585 = {1{`RANDOM}};
  _T_1981_re = _RAND_3585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3586 = {1{`RANDOM}};
  _T_1981_im = _RAND_3586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3587 = {1{`RANDOM}};
  _T_1982_re = _RAND_3587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3588 = {1{`RANDOM}};
  _T_1982_im = _RAND_3588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3589 = {1{`RANDOM}};
  _T_1983_re = _RAND_3589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3590 = {1{`RANDOM}};
  _T_1983_im = _RAND_3590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3591 = {1{`RANDOM}};
  _T_1984_re = _RAND_3591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3592 = {1{`RANDOM}};
  _T_1984_im = _RAND_3592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3593 = {1{`RANDOM}};
  _T_1985_re = _RAND_3593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3594 = {1{`RANDOM}};
  _T_1985_im = _RAND_3594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3595 = {1{`RANDOM}};
  _T_1986_re = _RAND_3595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3596 = {1{`RANDOM}};
  _T_1986_im = _RAND_3596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3597 = {1{`RANDOM}};
  _T_1987_re = _RAND_3597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3598 = {1{`RANDOM}};
  _T_1987_im = _RAND_3598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3599 = {1{`RANDOM}};
  _T_1988_re = _RAND_3599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3600 = {1{`RANDOM}};
  _T_1988_im = _RAND_3600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3601 = {1{`RANDOM}};
  _T_1989_re = _RAND_3601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3602 = {1{`RANDOM}};
  _T_1989_im = _RAND_3602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3603 = {1{`RANDOM}};
  _T_1990_re = _RAND_3603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3604 = {1{`RANDOM}};
  _T_1990_im = _RAND_3604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3605 = {1{`RANDOM}};
  _T_1991_re = _RAND_3605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3606 = {1{`RANDOM}};
  _T_1991_im = _RAND_3606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3607 = {1{`RANDOM}};
  _T_1992_re = _RAND_3607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3608 = {1{`RANDOM}};
  _T_1992_im = _RAND_3608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3609 = {1{`RANDOM}};
  _T_1993_re = _RAND_3609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3610 = {1{`RANDOM}};
  _T_1993_im = _RAND_3610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3611 = {1{`RANDOM}};
  _T_1994_re = _RAND_3611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3612 = {1{`RANDOM}};
  _T_1994_im = _RAND_3612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3613 = {1{`RANDOM}};
  _T_1995_re = _RAND_3613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3614 = {1{`RANDOM}};
  _T_1995_im = _RAND_3614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3615 = {1{`RANDOM}};
  _T_1996_re = _RAND_3615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3616 = {1{`RANDOM}};
  _T_1996_im = _RAND_3616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3617 = {1{`RANDOM}};
  _T_1997_re = _RAND_3617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3618 = {1{`RANDOM}};
  _T_1997_im = _RAND_3618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3619 = {1{`RANDOM}};
  _T_1998_re = _RAND_3619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3620 = {1{`RANDOM}};
  _T_1998_im = _RAND_3620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3621 = {1{`RANDOM}};
  _T_1999_re = _RAND_3621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3622 = {1{`RANDOM}};
  _T_1999_im = _RAND_3622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3623 = {1{`RANDOM}};
  _T_2000_re = _RAND_3623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3624 = {1{`RANDOM}};
  _T_2000_im = _RAND_3624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3625 = {1{`RANDOM}};
  _T_2001_re = _RAND_3625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3626 = {1{`RANDOM}};
  _T_2001_im = _RAND_3626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3627 = {1{`RANDOM}};
  _T_2002_re = _RAND_3627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3628 = {1{`RANDOM}};
  _T_2002_im = _RAND_3628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3629 = {1{`RANDOM}};
  _T_2003_re = _RAND_3629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3630 = {1{`RANDOM}};
  _T_2003_im = _RAND_3630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3631 = {1{`RANDOM}};
  _T_2004_re = _RAND_3631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3632 = {1{`RANDOM}};
  _T_2004_im = _RAND_3632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3633 = {1{`RANDOM}};
  _T_2005_re = _RAND_3633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3634 = {1{`RANDOM}};
  _T_2005_im = _RAND_3634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3635 = {1{`RANDOM}};
  _T_2006_re = _RAND_3635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3636 = {1{`RANDOM}};
  _T_2006_im = _RAND_3636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3637 = {1{`RANDOM}};
  _T_2007_re = _RAND_3637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3638 = {1{`RANDOM}};
  _T_2007_im = _RAND_3638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3639 = {1{`RANDOM}};
  _T_2008_re = _RAND_3639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3640 = {1{`RANDOM}};
  _T_2008_im = _RAND_3640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3641 = {1{`RANDOM}};
  _T_2009_re = _RAND_3641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3642 = {1{`RANDOM}};
  _T_2009_im = _RAND_3642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3643 = {1{`RANDOM}};
  _T_2010_re = _RAND_3643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3644 = {1{`RANDOM}};
  _T_2010_im = _RAND_3644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3645 = {1{`RANDOM}};
  _T_2011_re = _RAND_3645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3646 = {1{`RANDOM}};
  _T_2011_im = _RAND_3646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3647 = {1{`RANDOM}};
  _T_2012_re = _RAND_3647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3648 = {1{`RANDOM}};
  _T_2012_im = _RAND_3648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3649 = {1{`RANDOM}};
  _T_2013_re = _RAND_3649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3650 = {1{`RANDOM}};
  _T_2013_im = _RAND_3650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3651 = {1{`RANDOM}};
  _T_2014_re = _RAND_3651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3652 = {1{`RANDOM}};
  _T_2014_im = _RAND_3652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3653 = {1{`RANDOM}};
  _T_2015_re = _RAND_3653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3654 = {1{`RANDOM}};
  _T_2015_im = _RAND_3654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3655 = {1{`RANDOM}};
  _T_2016_re = _RAND_3655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3656 = {1{`RANDOM}};
  _T_2016_im = _RAND_3656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3657 = {1{`RANDOM}};
  _T_2017_re = _RAND_3657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3658 = {1{`RANDOM}};
  _T_2017_im = _RAND_3658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3659 = {1{`RANDOM}};
  _T_2018_re = _RAND_3659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3660 = {1{`RANDOM}};
  _T_2018_im = _RAND_3660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3661 = {1{`RANDOM}};
  _T_2019_re = _RAND_3661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3662 = {1{`RANDOM}};
  _T_2019_im = _RAND_3662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3663 = {1{`RANDOM}};
  _T_2020_re = _RAND_3663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3664 = {1{`RANDOM}};
  _T_2020_im = _RAND_3664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3665 = {1{`RANDOM}};
  _T_2021_re = _RAND_3665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3666 = {1{`RANDOM}};
  _T_2021_im = _RAND_3666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3667 = {1{`RANDOM}};
  _T_2022_re = _RAND_3667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3668 = {1{`RANDOM}};
  _T_2022_im = _RAND_3668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3669 = {1{`RANDOM}};
  _T_2023_re = _RAND_3669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3670 = {1{`RANDOM}};
  _T_2023_im = _RAND_3670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3671 = {1{`RANDOM}};
  _T_2024_re = _RAND_3671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3672 = {1{`RANDOM}};
  _T_2024_im = _RAND_3672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3673 = {1{`RANDOM}};
  _T_2025_re = _RAND_3673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3674 = {1{`RANDOM}};
  _T_2025_im = _RAND_3674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3675 = {1{`RANDOM}};
  _T_2026_re = _RAND_3675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3676 = {1{`RANDOM}};
  _T_2026_im = _RAND_3676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3677 = {1{`RANDOM}};
  _T_2027_re = _RAND_3677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3678 = {1{`RANDOM}};
  _T_2027_im = _RAND_3678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3679 = {1{`RANDOM}};
  _T_2028_re = _RAND_3679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3680 = {1{`RANDOM}};
  _T_2028_im = _RAND_3680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3681 = {1{`RANDOM}};
  _T_2029_re = _RAND_3681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3682 = {1{`RANDOM}};
  _T_2029_im = _RAND_3682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3683 = {1{`RANDOM}};
  _T_2030_re = _RAND_3683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3684 = {1{`RANDOM}};
  _T_2030_im = _RAND_3684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3685 = {1{`RANDOM}};
  _T_2031_re = _RAND_3685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3686 = {1{`RANDOM}};
  _T_2031_im = _RAND_3686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3687 = {1{`RANDOM}};
  _T_2032_re = _RAND_3687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3688 = {1{`RANDOM}};
  _T_2032_im = _RAND_3688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3689 = {1{`RANDOM}};
  _T_2033_re = _RAND_3689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3690 = {1{`RANDOM}};
  _T_2033_im = _RAND_3690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3691 = {1{`RANDOM}};
  _T_2034_re = _RAND_3691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3692 = {1{`RANDOM}};
  _T_2034_im = _RAND_3692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3693 = {1{`RANDOM}};
  _T_2035_re = _RAND_3693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3694 = {1{`RANDOM}};
  _T_2035_im = _RAND_3694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3695 = {1{`RANDOM}};
  _T_2036_re = _RAND_3695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3696 = {1{`RANDOM}};
  _T_2036_im = _RAND_3696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3697 = {1{`RANDOM}};
  _T_2037_re = _RAND_3697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3698 = {1{`RANDOM}};
  _T_2037_im = _RAND_3698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3699 = {1{`RANDOM}};
  _T_2038_re = _RAND_3699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3700 = {1{`RANDOM}};
  _T_2038_im = _RAND_3700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3701 = {1{`RANDOM}};
  _T_2039_re = _RAND_3701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3702 = {1{`RANDOM}};
  _T_2039_im = _RAND_3702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3703 = {1{`RANDOM}};
  _T_2040_re = _RAND_3703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3704 = {1{`RANDOM}};
  _T_2040_im = _RAND_3704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3705 = {1{`RANDOM}};
  _T_2041_re = _RAND_3705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3706 = {1{`RANDOM}};
  _T_2041_im = _RAND_3706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3707 = {1{`RANDOM}};
  _T_2042_re = _RAND_3707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3708 = {1{`RANDOM}};
  _T_2042_im = _RAND_3708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3709 = {1{`RANDOM}};
  _T_2043_re = _RAND_3709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3710 = {1{`RANDOM}};
  _T_2043_im = _RAND_3710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3711 = {1{`RANDOM}};
  _T_2044_re = _RAND_3711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3712 = {1{`RANDOM}};
  _T_2044_im = _RAND_3712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3713 = {1{`RANDOM}};
  _T_2045_re = _RAND_3713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3714 = {1{`RANDOM}};
  _T_2045_im = _RAND_3714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3715 = {1{`RANDOM}};
  _T_2046_re = _RAND_3715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3716 = {1{`RANDOM}};
  _T_2046_im = _RAND_3716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3717 = {1{`RANDOM}};
  _T_2047_re = _RAND_3717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3718 = {1{`RANDOM}};
  _T_2047_im = _RAND_3718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3719 = {1{`RANDOM}};
  _T_2048_re = _RAND_3719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3720 = {1{`RANDOM}};
  _T_2048_im = _RAND_3720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3721 = {1{`RANDOM}};
  _T_2049_re = _RAND_3721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3722 = {1{`RANDOM}};
  _T_2049_im = _RAND_3722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3723 = {1{`RANDOM}};
  _T_2050_re = _RAND_3723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3724 = {1{`RANDOM}};
  _T_2050_im = _RAND_3724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3725 = {1{`RANDOM}};
  _T_2051_re = _RAND_3725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3726 = {1{`RANDOM}};
  _T_2051_im = _RAND_3726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3727 = {1{`RANDOM}};
  _T_2052_re = _RAND_3727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3728 = {1{`RANDOM}};
  _T_2052_im = _RAND_3728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3729 = {1{`RANDOM}};
  _T_2053_re = _RAND_3729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3730 = {1{`RANDOM}};
  _T_2053_im = _RAND_3730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3731 = {1{`RANDOM}};
  _T_2054_re = _RAND_3731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3732 = {1{`RANDOM}};
  _T_2054_im = _RAND_3732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3733 = {1{`RANDOM}};
  _T_2055_re = _RAND_3733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3734 = {1{`RANDOM}};
  _T_2055_im = _RAND_3734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3735 = {1{`RANDOM}};
  _T_2056_re = _RAND_3735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3736 = {1{`RANDOM}};
  _T_2056_im = _RAND_3736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3737 = {1{`RANDOM}};
  _T_2057_re = _RAND_3737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3738 = {1{`RANDOM}};
  _T_2057_im = _RAND_3738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3739 = {1{`RANDOM}};
  _T_2058_re = _RAND_3739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3740 = {1{`RANDOM}};
  _T_2058_im = _RAND_3740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3741 = {1{`RANDOM}};
  _T_2059_re = _RAND_3741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3742 = {1{`RANDOM}};
  _T_2059_im = _RAND_3742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3743 = {1{`RANDOM}};
  _T_2060_re = _RAND_3743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3744 = {1{`RANDOM}};
  _T_2060_im = _RAND_3744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3745 = {1{`RANDOM}};
  _T_2061_re = _RAND_3745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3746 = {1{`RANDOM}};
  _T_2061_im = _RAND_3746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3747 = {1{`RANDOM}};
  _T_2062_re = _RAND_3747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3748 = {1{`RANDOM}};
  _T_2062_im = _RAND_3748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3749 = {1{`RANDOM}};
  _T_2063_re = _RAND_3749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3750 = {1{`RANDOM}};
  _T_2063_im = _RAND_3750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3751 = {1{`RANDOM}};
  _T_2064_re = _RAND_3751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3752 = {1{`RANDOM}};
  _T_2064_im = _RAND_3752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3753 = {1{`RANDOM}};
  _T_2065_re = _RAND_3753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3754 = {1{`RANDOM}};
  _T_2065_im = _RAND_3754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3755 = {1{`RANDOM}};
  _T_2066_re = _RAND_3755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3756 = {1{`RANDOM}};
  _T_2066_im = _RAND_3756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3757 = {1{`RANDOM}};
  _T_2067_re = _RAND_3757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3758 = {1{`RANDOM}};
  _T_2067_im = _RAND_3758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3759 = {1{`RANDOM}};
  _T_2068_re = _RAND_3759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3760 = {1{`RANDOM}};
  _T_2068_im = _RAND_3760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3761 = {1{`RANDOM}};
  _T_2069_re = _RAND_3761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3762 = {1{`RANDOM}};
  _T_2069_im = _RAND_3762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3763 = {1{`RANDOM}};
  _T_2070_re = _RAND_3763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3764 = {1{`RANDOM}};
  _T_2070_im = _RAND_3764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3765 = {1{`RANDOM}};
  _T_2071_re = _RAND_3765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3766 = {1{`RANDOM}};
  _T_2071_im = _RAND_3766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3767 = {1{`RANDOM}};
  _T_2072_re = _RAND_3767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3768 = {1{`RANDOM}};
  _T_2072_im = _RAND_3768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3769 = {1{`RANDOM}};
  _T_2073_re = _RAND_3769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3770 = {1{`RANDOM}};
  _T_2073_im = _RAND_3770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3771 = {1{`RANDOM}};
  _T_2074_re = _RAND_3771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3772 = {1{`RANDOM}};
  _T_2074_im = _RAND_3772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3773 = {1{`RANDOM}};
  _T_2075_re = _RAND_3773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3774 = {1{`RANDOM}};
  _T_2075_im = _RAND_3774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3775 = {1{`RANDOM}};
  _T_2076_re = _RAND_3775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3776 = {1{`RANDOM}};
  _T_2076_im = _RAND_3776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3777 = {1{`RANDOM}};
  _T_2077_re = _RAND_3777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3778 = {1{`RANDOM}};
  _T_2077_im = _RAND_3778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3779 = {1{`RANDOM}};
  _T_2078_re = _RAND_3779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3780 = {1{`RANDOM}};
  _T_2078_im = _RAND_3780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3781 = {1{`RANDOM}};
  _T_2079_re = _RAND_3781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3782 = {1{`RANDOM}};
  _T_2079_im = _RAND_3782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3783 = {1{`RANDOM}};
  _T_2080_re = _RAND_3783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3784 = {1{`RANDOM}};
  _T_2080_im = _RAND_3784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3785 = {1{`RANDOM}};
  _T_2081_re = _RAND_3785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3786 = {1{`RANDOM}};
  _T_2081_im = _RAND_3786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3787 = {1{`RANDOM}};
  _T_2082_re = _RAND_3787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3788 = {1{`RANDOM}};
  _T_2082_im = _RAND_3788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3789 = {1{`RANDOM}};
  _T_2083_re = _RAND_3789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3790 = {1{`RANDOM}};
  _T_2083_im = _RAND_3790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3791 = {1{`RANDOM}};
  _T_2084_re = _RAND_3791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3792 = {1{`RANDOM}};
  _T_2084_im = _RAND_3792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3793 = {1{`RANDOM}};
  _T_2085_re = _RAND_3793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3794 = {1{`RANDOM}};
  _T_2085_im = _RAND_3794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3795 = {1{`RANDOM}};
  _T_2086_re = _RAND_3795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3796 = {1{`RANDOM}};
  _T_2086_im = _RAND_3796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3797 = {1{`RANDOM}};
  _T_2087_re = _RAND_3797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3798 = {1{`RANDOM}};
  _T_2087_im = _RAND_3798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3799 = {1{`RANDOM}};
  _T_2088_re = _RAND_3799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3800 = {1{`RANDOM}};
  _T_2088_im = _RAND_3800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3801 = {1{`RANDOM}};
  _T_2089_re = _RAND_3801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3802 = {1{`RANDOM}};
  _T_2089_im = _RAND_3802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3803 = {1{`RANDOM}};
  _T_2090_re = _RAND_3803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3804 = {1{`RANDOM}};
  _T_2090_im = _RAND_3804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3805 = {1{`RANDOM}};
  _T_2091_re = _RAND_3805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3806 = {1{`RANDOM}};
  _T_2091_im = _RAND_3806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3807 = {1{`RANDOM}};
  _T_2092_re = _RAND_3807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3808 = {1{`RANDOM}};
  _T_2092_im = _RAND_3808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3809 = {1{`RANDOM}};
  _T_2093_re = _RAND_3809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3810 = {1{`RANDOM}};
  _T_2093_im = _RAND_3810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3811 = {1{`RANDOM}};
  _T_2094_re = _RAND_3811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3812 = {1{`RANDOM}};
  _T_2094_im = _RAND_3812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3813 = {1{`RANDOM}};
  _T_2095_re = _RAND_3813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3814 = {1{`RANDOM}};
  _T_2095_im = _RAND_3814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3815 = {1{`RANDOM}};
  _T_2096_re = _RAND_3815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3816 = {1{`RANDOM}};
  _T_2096_im = _RAND_3816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3817 = {1{`RANDOM}};
  _T_2097_re = _RAND_3817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3818 = {1{`RANDOM}};
  _T_2097_im = _RAND_3818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3819 = {1{`RANDOM}};
  _T_2098_re = _RAND_3819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3820 = {1{`RANDOM}};
  _T_2098_im = _RAND_3820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3821 = {1{`RANDOM}};
  _T_2099_re = _RAND_3821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3822 = {1{`RANDOM}};
  _T_2099_im = _RAND_3822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3823 = {1{`RANDOM}};
  _T_2100_re = _RAND_3823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3824 = {1{`RANDOM}};
  _T_2100_im = _RAND_3824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3825 = {1{`RANDOM}};
  _T_2101_re = _RAND_3825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3826 = {1{`RANDOM}};
  _T_2101_im = _RAND_3826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3827 = {1{`RANDOM}};
  _T_2102_re = _RAND_3827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3828 = {1{`RANDOM}};
  _T_2102_im = _RAND_3828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3829 = {1{`RANDOM}};
  _T_2103_re = _RAND_3829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3830 = {1{`RANDOM}};
  _T_2103_im = _RAND_3830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3831 = {1{`RANDOM}};
  _T_2104_re = _RAND_3831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3832 = {1{`RANDOM}};
  _T_2104_im = _RAND_3832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3833 = {1{`RANDOM}};
  _T_2105_re = _RAND_3833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3834 = {1{`RANDOM}};
  _T_2105_im = _RAND_3834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3835 = {1{`RANDOM}};
  _T_2106_re = _RAND_3835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3836 = {1{`RANDOM}};
  _T_2106_im = _RAND_3836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3837 = {1{`RANDOM}};
  _T_2107_re = _RAND_3837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3838 = {1{`RANDOM}};
  _T_2107_im = _RAND_3838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3839 = {1{`RANDOM}};
  _T_2108_re = _RAND_3839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3840 = {1{`RANDOM}};
  _T_2108_im = _RAND_3840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3841 = {1{`RANDOM}};
  _T_2109_re = _RAND_3841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3842 = {1{`RANDOM}};
  _T_2109_im = _RAND_3842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3843 = {1{`RANDOM}};
  _T_2110_re = _RAND_3843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3844 = {1{`RANDOM}};
  _T_2110_im = _RAND_3844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3845 = {1{`RANDOM}};
  _T_2111_re = _RAND_3845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3846 = {1{`RANDOM}};
  _T_2111_im = _RAND_3846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3847 = {1{`RANDOM}};
  _T_2112_re = _RAND_3847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3848 = {1{`RANDOM}};
  _T_2112_im = _RAND_3848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3849 = {1{`RANDOM}};
  _T_2113_re = _RAND_3849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3850 = {1{`RANDOM}};
  _T_2113_im = _RAND_3850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3851 = {1{`RANDOM}};
  _T_2114_re = _RAND_3851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3852 = {1{`RANDOM}};
  _T_2114_im = _RAND_3852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3853 = {1{`RANDOM}};
  _T_2115_re = _RAND_3853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3854 = {1{`RANDOM}};
  _T_2115_im = _RAND_3854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3855 = {1{`RANDOM}};
  _T_2116_re = _RAND_3855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3856 = {1{`RANDOM}};
  _T_2116_im = _RAND_3856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3857 = {1{`RANDOM}};
  _T_2117_re = _RAND_3857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3858 = {1{`RANDOM}};
  _T_2117_im = _RAND_3858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3859 = {1{`RANDOM}};
  _T_2118_re = _RAND_3859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3860 = {1{`RANDOM}};
  _T_2118_im = _RAND_3860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3861 = {1{`RANDOM}};
  _T_2119_re = _RAND_3861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3862 = {1{`RANDOM}};
  _T_2119_im = _RAND_3862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3863 = {1{`RANDOM}};
  _T_2120_re = _RAND_3863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3864 = {1{`RANDOM}};
  _T_2120_im = _RAND_3864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3865 = {1{`RANDOM}};
  _T_2121_re = _RAND_3865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3866 = {1{`RANDOM}};
  _T_2121_im = _RAND_3866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3867 = {1{`RANDOM}};
  _T_2122_re = _RAND_3867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3868 = {1{`RANDOM}};
  _T_2122_im = _RAND_3868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3869 = {1{`RANDOM}};
  _T_2123_re = _RAND_3869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3870 = {1{`RANDOM}};
  _T_2123_im = _RAND_3870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3871 = {1{`RANDOM}};
  _T_2124_re = _RAND_3871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3872 = {1{`RANDOM}};
  _T_2124_im = _RAND_3872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3873 = {1{`RANDOM}};
  _T_2125_re = _RAND_3873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3874 = {1{`RANDOM}};
  _T_2125_im = _RAND_3874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3875 = {1{`RANDOM}};
  _T_2126_re = _RAND_3875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3876 = {1{`RANDOM}};
  _T_2126_im = _RAND_3876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3877 = {1{`RANDOM}};
  _T_2127_re = _RAND_3877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3878 = {1{`RANDOM}};
  _T_2127_im = _RAND_3878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3879 = {1{`RANDOM}};
  _T_2128_re = _RAND_3879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3880 = {1{`RANDOM}};
  _T_2128_im = _RAND_3880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3881 = {1{`RANDOM}};
  _T_2129_re = _RAND_3881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3882 = {1{`RANDOM}};
  _T_2129_im = _RAND_3882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3883 = {1{`RANDOM}};
  _T_2130_re = _RAND_3883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3884 = {1{`RANDOM}};
  _T_2130_im = _RAND_3884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3885 = {1{`RANDOM}};
  _T_2131_re = _RAND_3885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3886 = {1{`RANDOM}};
  _T_2131_im = _RAND_3886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3887 = {1{`RANDOM}};
  _T_2132_re = _RAND_3887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3888 = {1{`RANDOM}};
  _T_2132_im = _RAND_3888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3889 = {1{`RANDOM}};
  _T_2133_re = _RAND_3889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3890 = {1{`RANDOM}};
  _T_2133_im = _RAND_3890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3891 = {1{`RANDOM}};
  _T_2134_re = _RAND_3891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3892 = {1{`RANDOM}};
  _T_2134_im = _RAND_3892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3893 = {1{`RANDOM}};
  _T_2135_re = _RAND_3893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3894 = {1{`RANDOM}};
  _T_2135_im = _RAND_3894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3895 = {1{`RANDOM}};
  _T_2136_re = _RAND_3895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3896 = {1{`RANDOM}};
  _T_2136_im = _RAND_3896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3897 = {1{`RANDOM}};
  _T_2137_re = _RAND_3897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3898 = {1{`RANDOM}};
  _T_2137_im = _RAND_3898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3899 = {1{`RANDOM}};
  _T_2138_re = _RAND_3899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3900 = {1{`RANDOM}};
  _T_2138_im = _RAND_3900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3901 = {1{`RANDOM}};
  _T_2139_re = _RAND_3901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3902 = {1{`RANDOM}};
  _T_2139_im = _RAND_3902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3903 = {1{`RANDOM}};
  _T_2140_re = _RAND_3903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3904 = {1{`RANDOM}};
  _T_2140_im = _RAND_3904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3905 = {1{`RANDOM}};
  _T_2141_re = _RAND_3905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3906 = {1{`RANDOM}};
  _T_2141_im = _RAND_3906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3907 = {1{`RANDOM}};
  _T_2142_re = _RAND_3907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3908 = {1{`RANDOM}};
  _T_2142_im = _RAND_3908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3909 = {1{`RANDOM}};
  _T_2143_re = _RAND_3909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3910 = {1{`RANDOM}};
  _T_2143_im = _RAND_3910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3911 = {1{`RANDOM}};
  _T_2144_re = _RAND_3911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3912 = {1{`RANDOM}};
  _T_2144_im = _RAND_3912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3913 = {1{`RANDOM}};
  _T_2145_re = _RAND_3913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3914 = {1{`RANDOM}};
  _T_2145_im = _RAND_3914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3915 = {1{`RANDOM}};
  _T_2146_re = _RAND_3915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3916 = {1{`RANDOM}};
  _T_2146_im = _RAND_3916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3917 = {1{`RANDOM}};
  _T_2147_re = _RAND_3917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3918 = {1{`RANDOM}};
  _T_2147_im = _RAND_3918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3919 = {1{`RANDOM}};
  _T_2148_re = _RAND_3919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3920 = {1{`RANDOM}};
  _T_2148_im = _RAND_3920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3921 = {1{`RANDOM}};
  _T_2149_re = _RAND_3921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3922 = {1{`RANDOM}};
  _T_2149_im = _RAND_3922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3923 = {1{`RANDOM}};
  _T_2150_re = _RAND_3923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3924 = {1{`RANDOM}};
  _T_2150_im = _RAND_3924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3925 = {1{`RANDOM}};
  _T_2151_re = _RAND_3925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3926 = {1{`RANDOM}};
  _T_2151_im = _RAND_3926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3927 = {1{`RANDOM}};
  _T_2152_re = _RAND_3927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3928 = {1{`RANDOM}};
  _T_2152_im = _RAND_3928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3929 = {1{`RANDOM}};
  _T_2153_re = _RAND_3929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3930 = {1{`RANDOM}};
  _T_2153_im = _RAND_3930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3931 = {1{`RANDOM}};
  _T_2154_re = _RAND_3931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3932 = {1{`RANDOM}};
  _T_2154_im = _RAND_3932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3933 = {1{`RANDOM}};
  _T_2155_re = _RAND_3933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3934 = {1{`RANDOM}};
  _T_2155_im = _RAND_3934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3935 = {1{`RANDOM}};
  _T_2156_re = _RAND_3935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3936 = {1{`RANDOM}};
  _T_2156_im = _RAND_3936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3937 = {1{`RANDOM}};
  _T_2157_re = _RAND_3937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3938 = {1{`RANDOM}};
  _T_2157_im = _RAND_3938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3939 = {1{`RANDOM}};
  _T_2158_re = _RAND_3939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3940 = {1{`RANDOM}};
  _T_2158_im = _RAND_3940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3941 = {1{`RANDOM}};
  _T_2159_re = _RAND_3941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3942 = {1{`RANDOM}};
  _T_2159_im = _RAND_3942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3943 = {1{`RANDOM}};
  _T_2160_re = _RAND_3943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3944 = {1{`RANDOM}};
  _T_2160_im = _RAND_3944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3945 = {1{`RANDOM}};
  _T_2161_re = _RAND_3945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3946 = {1{`RANDOM}};
  _T_2161_im = _RAND_3946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3947 = {1{`RANDOM}};
  _T_2162_re = _RAND_3947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3948 = {1{`RANDOM}};
  _T_2162_im = _RAND_3948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3949 = {1{`RANDOM}};
  _T_2163_re = _RAND_3949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3950 = {1{`RANDOM}};
  _T_2163_im = _RAND_3950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3951 = {1{`RANDOM}};
  _T_2164_re = _RAND_3951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3952 = {1{`RANDOM}};
  _T_2164_im = _RAND_3952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3953 = {1{`RANDOM}};
  _T_2165_re = _RAND_3953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3954 = {1{`RANDOM}};
  _T_2165_im = _RAND_3954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3955 = {1{`RANDOM}};
  _T_2166_re = _RAND_3955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3956 = {1{`RANDOM}};
  _T_2166_im = _RAND_3956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3957 = {1{`RANDOM}};
  _T_2167_re = _RAND_3957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3958 = {1{`RANDOM}};
  _T_2167_im = _RAND_3958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3959 = {1{`RANDOM}};
  _T_2168_re = _RAND_3959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3960 = {1{`RANDOM}};
  _T_2168_im = _RAND_3960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3961 = {1{`RANDOM}};
  _T_2169_re = _RAND_3961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3962 = {1{`RANDOM}};
  _T_2169_im = _RAND_3962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3963 = {1{`RANDOM}};
  _T_2170_re = _RAND_3963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3964 = {1{`RANDOM}};
  _T_2170_im = _RAND_3964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3965 = {1{`RANDOM}};
  _T_2171_re = _RAND_3965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3966 = {1{`RANDOM}};
  _T_2171_im = _RAND_3966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3967 = {1{`RANDOM}};
  _T_2172_re = _RAND_3967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3968 = {1{`RANDOM}};
  _T_2172_im = _RAND_3968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3969 = {1{`RANDOM}};
  _T_2173_re = _RAND_3969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3970 = {1{`RANDOM}};
  _T_2173_im = _RAND_3970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3971 = {1{`RANDOM}};
  _T_2174_re = _RAND_3971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3972 = {1{`RANDOM}};
  _T_2174_im = _RAND_3972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3973 = {1{`RANDOM}};
  _T_2175_re = _RAND_3973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3974 = {1{`RANDOM}};
  _T_2175_im = _RAND_3974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3975 = {1{`RANDOM}};
  _T_2176_re = _RAND_3975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3976 = {1{`RANDOM}};
  _T_2176_im = _RAND_3976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3977 = {1{`RANDOM}};
  _T_2177_re = _RAND_3977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3978 = {1{`RANDOM}};
  _T_2177_im = _RAND_3978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3979 = {1{`RANDOM}};
  _T_2178_re = _RAND_3979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3980 = {1{`RANDOM}};
  _T_2178_im = _RAND_3980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3981 = {1{`RANDOM}};
  _T_2179_re = _RAND_3981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3982 = {1{`RANDOM}};
  _T_2179_im = _RAND_3982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3983 = {1{`RANDOM}};
  _T_2180_re = _RAND_3983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3984 = {1{`RANDOM}};
  _T_2180_im = _RAND_3984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3985 = {1{`RANDOM}};
  _T_2181_re = _RAND_3985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3986 = {1{`RANDOM}};
  _T_2181_im = _RAND_3986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3987 = {1{`RANDOM}};
  _T_2182_re = _RAND_3987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3988 = {1{`RANDOM}};
  _T_2182_im = _RAND_3988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3989 = {1{`RANDOM}};
  _T_2183_re = _RAND_3989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3990 = {1{`RANDOM}};
  _T_2183_im = _RAND_3990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3991 = {1{`RANDOM}};
  _T_2184_re = _RAND_3991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3992 = {1{`RANDOM}};
  _T_2184_im = _RAND_3992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3993 = {1{`RANDOM}};
  _T_2185_re = _RAND_3993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3994 = {1{`RANDOM}};
  _T_2185_im = _RAND_3994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3995 = {1{`RANDOM}};
  _T_2186_re = _RAND_3995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3996 = {1{`RANDOM}};
  _T_2186_im = _RAND_3996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3997 = {1{`RANDOM}};
  _T_2187_re = _RAND_3997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3998 = {1{`RANDOM}};
  _T_2187_im = _RAND_3998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3999 = {1{`RANDOM}};
  _T_2188_re = _RAND_3999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4000 = {1{`RANDOM}};
  _T_2188_im = _RAND_4000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4001 = {1{`RANDOM}};
  _T_2189_re = _RAND_4001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4002 = {1{`RANDOM}};
  _T_2189_im = _RAND_4002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4003 = {1{`RANDOM}};
  _T_2190_re = _RAND_4003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4004 = {1{`RANDOM}};
  _T_2190_im = _RAND_4004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4005 = {1{`RANDOM}};
  _T_2191_re = _RAND_4005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4006 = {1{`RANDOM}};
  _T_2191_im = _RAND_4006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4007 = {1{`RANDOM}};
  _T_2192_re = _RAND_4007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4008 = {1{`RANDOM}};
  _T_2192_im = _RAND_4008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4009 = {1{`RANDOM}};
  _T_2193_re = _RAND_4009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4010 = {1{`RANDOM}};
  _T_2193_im = _RAND_4010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4011 = {1{`RANDOM}};
  _T_2194_re = _RAND_4011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4012 = {1{`RANDOM}};
  _T_2194_im = _RAND_4012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4013 = {1{`RANDOM}};
  _T_2195_re = _RAND_4013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4014 = {1{`RANDOM}};
  _T_2195_im = _RAND_4014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4015 = {1{`RANDOM}};
  _T_2196_re = _RAND_4015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4016 = {1{`RANDOM}};
  _T_2196_im = _RAND_4016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4017 = {1{`RANDOM}};
  _T_2197_re = _RAND_4017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4018 = {1{`RANDOM}};
  _T_2197_im = _RAND_4018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4019 = {1{`RANDOM}};
  _T_2198_re = _RAND_4019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4020 = {1{`RANDOM}};
  _T_2198_im = _RAND_4020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4021 = {1{`RANDOM}};
  _T_2199_re = _RAND_4021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4022 = {1{`RANDOM}};
  _T_2199_im = _RAND_4022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4023 = {1{`RANDOM}};
  _T_2200_re = _RAND_4023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4024 = {1{`RANDOM}};
  _T_2200_im = _RAND_4024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4025 = {1{`RANDOM}};
  _T_2201_re = _RAND_4025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4026 = {1{`RANDOM}};
  _T_2201_im = _RAND_4026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4027 = {1{`RANDOM}};
  _T_2202_re = _RAND_4027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4028 = {1{`RANDOM}};
  _T_2202_im = _RAND_4028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4029 = {1{`RANDOM}};
  _T_2203_re = _RAND_4029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4030 = {1{`RANDOM}};
  _T_2203_im = _RAND_4030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4031 = {1{`RANDOM}};
  _T_2204_re = _RAND_4031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4032 = {1{`RANDOM}};
  _T_2204_im = _RAND_4032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4033 = {1{`RANDOM}};
  _T_2205_re = _RAND_4033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4034 = {1{`RANDOM}};
  _T_2205_im = _RAND_4034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4035 = {1{`RANDOM}};
  _T_2206_re = _RAND_4035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4036 = {1{`RANDOM}};
  _T_2206_im = _RAND_4036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4037 = {1{`RANDOM}};
  _T_2207_re = _RAND_4037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4038 = {1{`RANDOM}};
  _T_2207_im = _RAND_4038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4039 = {1{`RANDOM}};
  _T_2208_re = _RAND_4039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4040 = {1{`RANDOM}};
  _T_2208_im = _RAND_4040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4041 = {1{`RANDOM}};
  _T_2209_re = _RAND_4041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4042 = {1{`RANDOM}};
  _T_2209_im = _RAND_4042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4043 = {1{`RANDOM}};
  _T_2210_re = _RAND_4043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4044 = {1{`RANDOM}};
  _T_2210_im = _RAND_4044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4045 = {1{`RANDOM}};
  _T_2211_re = _RAND_4045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4046 = {1{`RANDOM}};
  _T_2211_im = _RAND_4046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4047 = {1{`RANDOM}};
  _T_2212_re = _RAND_4047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4048 = {1{`RANDOM}};
  _T_2212_im = _RAND_4048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4049 = {1{`RANDOM}};
  _T_2213_re = _RAND_4049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4050 = {1{`RANDOM}};
  _T_2213_im = _RAND_4050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4051 = {1{`RANDOM}};
  _T_2214_re = _RAND_4051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4052 = {1{`RANDOM}};
  _T_2214_im = _RAND_4052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4053 = {1{`RANDOM}};
  _T_2215_re = _RAND_4053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4054 = {1{`RANDOM}};
  _T_2215_im = _RAND_4054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4055 = {1{`RANDOM}};
  _T_2216_re = _RAND_4055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4056 = {1{`RANDOM}};
  _T_2216_im = _RAND_4056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4057 = {1{`RANDOM}};
  _T_2217_re = _RAND_4057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4058 = {1{`RANDOM}};
  _T_2217_im = _RAND_4058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4059 = {1{`RANDOM}};
  _T_2218_re = _RAND_4059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4060 = {1{`RANDOM}};
  _T_2218_im = _RAND_4060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4061 = {1{`RANDOM}};
  _T_2219_re = _RAND_4061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4062 = {1{`RANDOM}};
  _T_2219_im = _RAND_4062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4063 = {1{`RANDOM}};
  _T_2220_re = _RAND_4063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4064 = {1{`RANDOM}};
  _T_2220_im = _RAND_4064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4065 = {1{`RANDOM}};
  _T_2221_re = _RAND_4065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4066 = {1{`RANDOM}};
  _T_2221_im = _RAND_4066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4067 = {1{`RANDOM}};
  _T_2222_re = _RAND_4067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4068 = {1{`RANDOM}};
  _T_2222_im = _RAND_4068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4069 = {1{`RANDOM}};
  _T_2223_re = _RAND_4069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4070 = {1{`RANDOM}};
  _T_2223_im = _RAND_4070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4071 = {1{`RANDOM}};
  _T_2224_re = _RAND_4071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4072 = {1{`RANDOM}};
  _T_2224_im = _RAND_4072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4073 = {1{`RANDOM}};
  _T_2225_re = _RAND_4073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4074 = {1{`RANDOM}};
  _T_2225_im = _RAND_4074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4075 = {1{`RANDOM}};
  _T_2226_re = _RAND_4075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4076 = {1{`RANDOM}};
  _T_2226_im = _RAND_4076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4077 = {1{`RANDOM}};
  _T_2227_re = _RAND_4077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4078 = {1{`RANDOM}};
  _T_2227_im = _RAND_4078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4079 = {1{`RANDOM}};
  _T_2228_re = _RAND_4079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4080 = {1{`RANDOM}};
  _T_2228_im = _RAND_4080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4081 = {1{`RANDOM}};
  _T_2229_re = _RAND_4081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4082 = {1{`RANDOM}};
  _T_2229_im = _RAND_4082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4083 = {1{`RANDOM}};
  _T_2230_re = _RAND_4083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4084 = {1{`RANDOM}};
  _T_2230_im = _RAND_4084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4085 = {1{`RANDOM}};
  _T_2231_re = _RAND_4085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4086 = {1{`RANDOM}};
  _T_2231_im = _RAND_4086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4087 = {1{`RANDOM}};
  _T_2232_re = _RAND_4087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4088 = {1{`RANDOM}};
  _T_2232_im = _RAND_4088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4089 = {1{`RANDOM}};
  _T_2233_re = _RAND_4089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4090 = {1{`RANDOM}};
  _T_2233_im = _RAND_4090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4091 = {1{`RANDOM}};
  _T_2234_re = _RAND_4091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4092 = {1{`RANDOM}};
  _T_2234_im = _RAND_4092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4093 = {1{`RANDOM}};
  _T_2235_re = _RAND_4093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4094 = {1{`RANDOM}};
  _T_2235_im = _RAND_4094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4095 = {1{`RANDOM}};
  _T_2236_re = _RAND_4095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4096 = {1{`RANDOM}};
  _T_2236_im = _RAND_4096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4097 = {1{`RANDOM}};
  _T_2237_re = _RAND_4097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4098 = {1{`RANDOM}};
  _T_2237_im = _RAND_4098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4099 = {1{`RANDOM}};
  _T_2238_re = _RAND_4099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4100 = {1{`RANDOM}};
  _T_2238_im = _RAND_4100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4101 = {1{`RANDOM}};
  _T_2239_re = _RAND_4101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4102 = {1{`RANDOM}};
  _T_2239_im = _RAND_4102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4103 = {1{`RANDOM}};
  _T_2242_re = _RAND_4103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4104 = {1{`RANDOM}};
  _T_2242_im = _RAND_4104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4105 = {1{`RANDOM}};
  _T_2243_re = _RAND_4105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4106 = {1{`RANDOM}};
  _T_2243_im = _RAND_4106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4107 = {1{`RANDOM}};
  _T_2244_re = _RAND_4107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4108 = {1{`RANDOM}};
  _T_2244_im = _RAND_4108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4109 = {1{`RANDOM}};
  _T_2245_re = _RAND_4109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4110 = {1{`RANDOM}};
  _T_2245_im = _RAND_4110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4111 = {1{`RANDOM}};
  _T_2246_re = _RAND_4111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4112 = {1{`RANDOM}};
  _T_2246_im = _RAND_4112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4113 = {1{`RANDOM}};
  _T_2247_re = _RAND_4113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4114 = {1{`RANDOM}};
  _T_2247_im = _RAND_4114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4115 = {1{`RANDOM}};
  _T_2248_re = _RAND_4115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4116 = {1{`RANDOM}};
  _T_2248_im = _RAND_4116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4117 = {1{`RANDOM}};
  _T_2249_re = _RAND_4117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4118 = {1{`RANDOM}};
  _T_2249_im = _RAND_4118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4119 = {1{`RANDOM}};
  _T_2250_re = _RAND_4119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4120 = {1{`RANDOM}};
  _T_2250_im = _RAND_4120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4121 = {1{`RANDOM}};
  _T_2251_re = _RAND_4121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4122 = {1{`RANDOM}};
  _T_2251_im = _RAND_4122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4123 = {1{`RANDOM}};
  _T_2252_re = _RAND_4123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4124 = {1{`RANDOM}};
  _T_2252_im = _RAND_4124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4125 = {1{`RANDOM}};
  _T_2253_re = _RAND_4125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4126 = {1{`RANDOM}};
  _T_2253_im = _RAND_4126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4127 = {1{`RANDOM}};
  _T_2254_re = _RAND_4127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4128 = {1{`RANDOM}};
  _T_2254_im = _RAND_4128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4129 = {1{`RANDOM}};
  _T_2255_re = _RAND_4129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4130 = {1{`RANDOM}};
  _T_2255_im = _RAND_4130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4131 = {1{`RANDOM}};
  _T_2256_re = _RAND_4131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4132 = {1{`RANDOM}};
  _T_2256_im = _RAND_4132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4133 = {1{`RANDOM}};
  _T_2257_re = _RAND_4133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4134 = {1{`RANDOM}};
  _T_2257_im = _RAND_4134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4135 = {1{`RANDOM}};
  _T_2258_re = _RAND_4135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4136 = {1{`RANDOM}};
  _T_2258_im = _RAND_4136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4137 = {1{`RANDOM}};
  _T_2259_re = _RAND_4137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4138 = {1{`RANDOM}};
  _T_2259_im = _RAND_4138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4139 = {1{`RANDOM}};
  _T_2260_re = _RAND_4139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4140 = {1{`RANDOM}};
  _T_2260_im = _RAND_4140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4141 = {1{`RANDOM}};
  _T_2261_re = _RAND_4141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4142 = {1{`RANDOM}};
  _T_2261_im = _RAND_4142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4143 = {1{`RANDOM}};
  _T_2262_re = _RAND_4143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4144 = {1{`RANDOM}};
  _T_2262_im = _RAND_4144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4145 = {1{`RANDOM}};
  _T_2263_re = _RAND_4145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4146 = {1{`RANDOM}};
  _T_2263_im = _RAND_4146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4147 = {1{`RANDOM}};
  _T_2264_re = _RAND_4147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4148 = {1{`RANDOM}};
  _T_2264_im = _RAND_4148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4149 = {1{`RANDOM}};
  _T_2265_re = _RAND_4149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4150 = {1{`RANDOM}};
  _T_2265_im = _RAND_4150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4151 = {1{`RANDOM}};
  _T_2266_re = _RAND_4151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4152 = {1{`RANDOM}};
  _T_2266_im = _RAND_4152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4153 = {1{`RANDOM}};
  _T_2267_re = _RAND_4153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4154 = {1{`RANDOM}};
  _T_2267_im = _RAND_4154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4155 = {1{`RANDOM}};
  _T_2268_re = _RAND_4155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4156 = {1{`RANDOM}};
  _T_2268_im = _RAND_4156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4157 = {1{`RANDOM}};
  _T_2269_re = _RAND_4157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4158 = {1{`RANDOM}};
  _T_2269_im = _RAND_4158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4159 = {1{`RANDOM}};
  _T_2270_re = _RAND_4159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4160 = {1{`RANDOM}};
  _T_2270_im = _RAND_4160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4161 = {1{`RANDOM}};
  _T_2271_re = _RAND_4161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4162 = {1{`RANDOM}};
  _T_2271_im = _RAND_4162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4163 = {1{`RANDOM}};
  _T_2272_re = _RAND_4163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4164 = {1{`RANDOM}};
  _T_2272_im = _RAND_4164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4165 = {1{`RANDOM}};
  _T_2273_re = _RAND_4165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4166 = {1{`RANDOM}};
  _T_2273_im = _RAND_4166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4167 = {1{`RANDOM}};
  _T_2274_re = _RAND_4167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4168 = {1{`RANDOM}};
  _T_2274_im = _RAND_4168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4169 = {1{`RANDOM}};
  _T_2275_re = _RAND_4169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4170 = {1{`RANDOM}};
  _T_2275_im = _RAND_4170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4171 = {1{`RANDOM}};
  _T_2276_re = _RAND_4171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4172 = {1{`RANDOM}};
  _T_2276_im = _RAND_4172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4173 = {1{`RANDOM}};
  _T_2277_re = _RAND_4173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4174 = {1{`RANDOM}};
  _T_2277_im = _RAND_4174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4175 = {1{`RANDOM}};
  _T_2278_re = _RAND_4175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4176 = {1{`RANDOM}};
  _T_2278_im = _RAND_4176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4177 = {1{`RANDOM}};
  _T_2279_re = _RAND_4177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4178 = {1{`RANDOM}};
  _T_2279_im = _RAND_4178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4179 = {1{`RANDOM}};
  _T_2280_re = _RAND_4179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4180 = {1{`RANDOM}};
  _T_2280_im = _RAND_4180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4181 = {1{`RANDOM}};
  _T_2281_re = _RAND_4181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4182 = {1{`RANDOM}};
  _T_2281_im = _RAND_4182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4183 = {1{`RANDOM}};
  _T_2282_re = _RAND_4183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4184 = {1{`RANDOM}};
  _T_2282_im = _RAND_4184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4185 = {1{`RANDOM}};
  _T_2283_re = _RAND_4185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4186 = {1{`RANDOM}};
  _T_2283_im = _RAND_4186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4187 = {1{`RANDOM}};
  _T_2284_re = _RAND_4187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4188 = {1{`RANDOM}};
  _T_2284_im = _RAND_4188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4189 = {1{`RANDOM}};
  _T_2285_re = _RAND_4189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4190 = {1{`RANDOM}};
  _T_2285_im = _RAND_4190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4191 = {1{`RANDOM}};
  _T_2286_re = _RAND_4191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4192 = {1{`RANDOM}};
  _T_2286_im = _RAND_4192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4193 = {1{`RANDOM}};
  _T_2287_re = _RAND_4193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4194 = {1{`RANDOM}};
  _T_2287_im = _RAND_4194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4195 = {1{`RANDOM}};
  _T_2288_re = _RAND_4195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4196 = {1{`RANDOM}};
  _T_2288_im = _RAND_4196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4197 = {1{`RANDOM}};
  _T_2289_re = _RAND_4197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4198 = {1{`RANDOM}};
  _T_2289_im = _RAND_4198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4199 = {1{`RANDOM}};
  _T_2290_re = _RAND_4199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4200 = {1{`RANDOM}};
  _T_2290_im = _RAND_4200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4201 = {1{`RANDOM}};
  _T_2291_re = _RAND_4201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4202 = {1{`RANDOM}};
  _T_2291_im = _RAND_4202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4203 = {1{`RANDOM}};
  _T_2292_re = _RAND_4203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4204 = {1{`RANDOM}};
  _T_2292_im = _RAND_4204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4205 = {1{`RANDOM}};
  _T_2293_re = _RAND_4205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4206 = {1{`RANDOM}};
  _T_2293_im = _RAND_4206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4207 = {1{`RANDOM}};
  _T_2294_re = _RAND_4207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4208 = {1{`RANDOM}};
  _T_2294_im = _RAND_4208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4209 = {1{`RANDOM}};
  _T_2295_re = _RAND_4209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4210 = {1{`RANDOM}};
  _T_2295_im = _RAND_4210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4211 = {1{`RANDOM}};
  _T_2296_re = _RAND_4211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4212 = {1{`RANDOM}};
  _T_2296_im = _RAND_4212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4213 = {1{`RANDOM}};
  _T_2297_re = _RAND_4213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4214 = {1{`RANDOM}};
  _T_2297_im = _RAND_4214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4215 = {1{`RANDOM}};
  _T_2298_re = _RAND_4215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4216 = {1{`RANDOM}};
  _T_2298_im = _RAND_4216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4217 = {1{`RANDOM}};
  _T_2299_re = _RAND_4217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4218 = {1{`RANDOM}};
  _T_2299_im = _RAND_4218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4219 = {1{`RANDOM}};
  _T_2300_re = _RAND_4219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4220 = {1{`RANDOM}};
  _T_2300_im = _RAND_4220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4221 = {1{`RANDOM}};
  _T_2301_re = _RAND_4221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4222 = {1{`RANDOM}};
  _T_2301_im = _RAND_4222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4223 = {1{`RANDOM}};
  _T_2302_re = _RAND_4223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4224 = {1{`RANDOM}};
  _T_2302_im = _RAND_4224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4225 = {1{`RANDOM}};
  _T_2303_re = _RAND_4225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4226 = {1{`RANDOM}};
  _T_2303_im = _RAND_4226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4227 = {1{`RANDOM}};
  _T_2304_re = _RAND_4227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4228 = {1{`RANDOM}};
  _T_2304_im = _RAND_4228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4229 = {1{`RANDOM}};
  _T_2305_re = _RAND_4229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4230 = {1{`RANDOM}};
  _T_2305_im = _RAND_4230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4231 = {1{`RANDOM}};
  _T_2306_re = _RAND_4231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4232 = {1{`RANDOM}};
  _T_2306_im = _RAND_4232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4233 = {1{`RANDOM}};
  _T_2307_re = _RAND_4233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4234 = {1{`RANDOM}};
  _T_2307_im = _RAND_4234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4235 = {1{`RANDOM}};
  _T_2308_re = _RAND_4235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4236 = {1{`RANDOM}};
  _T_2308_im = _RAND_4236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4237 = {1{`RANDOM}};
  _T_2309_re = _RAND_4237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4238 = {1{`RANDOM}};
  _T_2309_im = _RAND_4238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4239 = {1{`RANDOM}};
  _T_2310_re = _RAND_4239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4240 = {1{`RANDOM}};
  _T_2310_im = _RAND_4240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4241 = {1{`RANDOM}};
  _T_2311_re = _RAND_4241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4242 = {1{`RANDOM}};
  _T_2311_im = _RAND_4242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4243 = {1{`RANDOM}};
  _T_2312_re = _RAND_4243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4244 = {1{`RANDOM}};
  _T_2312_im = _RAND_4244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4245 = {1{`RANDOM}};
  _T_2313_re = _RAND_4245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4246 = {1{`RANDOM}};
  _T_2313_im = _RAND_4246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4247 = {1{`RANDOM}};
  _T_2314_re = _RAND_4247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4248 = {1{`RANDOM}};
  _T_2314_im = _RAND_4248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4249 = {1{`RANDOM}};
  _T_2315_re = _RAND_4249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4250 = {1{`RANDOM}};
  _T_2315_im = _RAND_4250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4251 = {1{`RANDOM}};
  _T_2316_re = _RAND_4251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4252 = {1{`RANDOM}};
  _T_2316_im = _RAND_4252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4253 = {1{`RANDOM}};
  _T_2317_re = _RAND_4253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4254 = {1{`RANDOM}};
  _T_2317_im = _RAND_4254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4255 = {1{`RANDOM}};
  _T_2318_re = _RAND_4255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4256 = {1{`RANDOM}};
  _T_2318_im = _RAND_4256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4257 = {1{`RANDOM}};
  _T_2319_re = _RAND_4257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4258 = {1{`RANDOM}};
  _T_2319_im = _RAND_4258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4259 = {1{`RANDOM}};
  _T_2320_re = _RAND_4259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4260 = {1{`RANDOM}};
  _T_2320_im = _RAND_4260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4261 = {1{`RANDOM}};
  _T_2321_re = _RAND_4261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4262 = {1{`RANDOM}};
  _T_2321_im = _RAND_4262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4263 = {1{`RANDOM}};
  _T_2322_re = _RAND_4263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4264 = {1{`RANDOM}};
  _T_2322_im = _RAND_4264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4265 = {1{`RANDOM}};
  _T_2323_re = _RAND_4265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4266 = {1{`RANDOM}};
  _T_2323_im = _RAND_4266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4267 = {1{`RANDOM}};
  _T_2324_re = _RAND_4267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4268 = {1{`RANDOM}};
  _T_2324_im = _RAND_4268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4269 = {1{`RANDOM}};
  _T_2325_re = _RAND_4269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4270 = {1{`RANDOM}};
  _T_2325_im = _RAND_4270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4271 = {1{`RANDOM}};
  _T_2326_re = _RAND_4271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4272 = {1{`RANDOM}};
  _T_2326_im = _RAND_4272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4273 = {1{`RANDOM}};
  _T_2327_re = _RAND_4273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4274 = {1{`RANDOM}};
  _T_2327_im = _RAND_4274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4275 = {1{`RANDOM}};
  _T_2328_re = _RAND_4275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4276 = {1{`RANDOM}};
  _T_2328_im = _RAND_4276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4277 = {1{`RANDOM}};
  _T_2329_re = _RAND_4277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4278 = {1{`RANDOM}};
  _T_2329_im = _RAND_4278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4279 = {1{`RANDOM}};
  _T_2330_re = _RAND_4279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4280 = {1{`RANDOM}};
  _T_2330_im = _RAND_4280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4281 = {1{`RANDOM}};
  _T_2331_re = _RAND_4281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4282 = {1{`RANDOM}};
  _T_2331_im = _RAND_4282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4283 = {1{`RANDOM}};
  _T_2332_re = _RAND_4283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4284 = {1{`RANDOM}};
  _T_2332_im = _RAND_4284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4285 = {1{`RANDOM}};
  _T_2333_re = _RAND_4285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4286 = {1{`RANDOM}};
  _T_2333_im = _RAND_4286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4287 = {1{`RANDOM}};
  _T_2334_re = _RAND_4287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4288 = {1{`RANDOM}};
  _T_2334_im = _RAND_4288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4289 = {1{`RANDOM}};
  _T_2335_re = _RAND_4289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4290 = {1{`RANDOM}};
  _T_2335_im = _RAND_4290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4291 = {1{`RANDOM}};
  _T_2336_re = _RAND_4291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4292 = {1{`RANDOM}};
  _T_2336_im = _RAND_4292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4293 = {1{`RANDOM}};
  _T_2337_re = _RAND_4293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4294 = {1{`RANDOM}};
  _T_2337_im = _RAND_4294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4295 = {1{`RANDOM}};
  _T_2338_re = _RAND_4295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4296 = {1{`RANDOM}};
  _T_2338_im = _RAND_4296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4297 = {1{`RANDOM}};
  _T_2339_re = _RAND_4297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4298 = {1{`RANDOM}};
  _T_2339_im = _RAND_4298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4299 = {1{`RANDOM}};
  _T_2340_re = _RAND_4299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4300 = {1{`RANDOM}};
  _T_2340_im = _RAND_4300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4301 = {1{`RANDOM}};
  _T_2341_re = _RAND_4301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4302 = {1{`RANDOM}};
  _T_2341_im = _RAND_4302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4303 = {1{`RANDOM}};
  _T_2342_re = _RAND_4303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4304 = {1{`RANDOM}};
  _T_2342_im = _RAND_4304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4305 = {1{`RANDOM}};
  _T_2343_re = _RAND_4305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4306 = {1{`RANDOM}};
  _T_2343_im = _RAND_4306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4307 = {1{`RANDOM}};
  _T_2344_re = _RAND_4307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4308 = {1{`RANDOM}};
  _T_2344_im = _RAND_4308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4309 = {1{`RANDOM}};
  _T_2345_re = _RAND_4309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4310 = {1{`RANDOM}};
  _T_2345_im = _RAND_4310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4311 = {1{`RANDOM}};
  _T_2346_re = _RAND_4311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4312 = {1{`RANDOM}};
  _T_2346_im = _RAND_4312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4313 = {1{`RANDOM}};
  _T_2347_re = _RAND_4313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4314 = {1{`RANDOM}};
  _T_2347_im = _RAND_4314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4315 = {1{`RANDOM}};
  _T_2348_re = _RAND_4315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4316 = {1{`RANDOM}};
  _T_2348_im = _RAND_4316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4317 = {1{`RANDOM}};
  _T_2349_re = _RAND_4317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4318 = {1{`RANDOM}};
  _T_2349_im = _RAND_4318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4319 = {1{`RANDOM}};
  _T_2350_re = _RAND_4319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4320 = {1{`RANDOM}};
  _T_2350_im = _RAND_4320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4321 = {1{`RANDOM}};
  _T_2351_re = _RAND_4321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4322 = {1{`RANDOM}};
  _T_2351_im = _RAND_4322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4323 = {1{`RANDOM}};
  _T_2352_re = _RAND_4323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4324 = {1{`RANDOM}};
  _T_2352_im = _RAND_4324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4325 = {1{`RANDOM}};
  _T_2353_re = _RAND_4325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4326 = {1{`RANDOM}};
  _T_2353_im = _RAND_4326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4327 = {1{`RANDOM}};
  _T_2354_re = _RAND_4327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4328 = {1{`RANDOM}};
  _T_2354_im = _RAND_4328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4329 = {1{`RANDOM}};
  _T_2355_re = _RAND_4329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4330 = {1{`RANDOM}};
  _T_2355_im = _RAND_4330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4331 = {1{`RANDOM}};
  _T_2356_re = _RAND_4331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4332 = {1{`RANDOM}};
  _T_2356_im = _RAND_4332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4333 = {1{`RANDOM}};
  _T_2357_re = _RAND_4333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4334 = {1{`RANDOM}};
  _T_2357_im = _RAND_4334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4335 = {1{`RANDOM}};
  _T_2358_re = _RAND_4335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4336 = {1{`RANDOM}};
  _T_2358_im = _RAND_4336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4337 = {1{`RANDOM}};
  _T_2359_re = _RAND_4337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4338 = {1{`RANDOM}};
  _T_2359_im = _RAND_4338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4339 = {1{`RANDOM}};
  _T_2360_re = _RAND_4339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4340 = {1{`RANDOM}};
  _T_2360_im = _RAND_4340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4341 = {1{`RANDOM}};
  _T_2361_re = _RAND_4341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4342 = {1{`RANDOM}};
  _T_2361_im = _RAND_4342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4343 = {1{`RANDOM}};
  _T_2362_re = _RAND_4343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4344 = {1{`RANDOM}};
  _T_2362_im = _RAND_4344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4345 = {1{`RANDOM}};
  _T_2363_re = _RAND_4345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4346 = {1{`RANDOM}};
  _T_2363_im = _RAND_4346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4347 = {1{`RANDOM}};
  _T_2364_re = _RAND_4347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4348 = {1{`RANDOM}};
  _T_2364_im = _RAND_4348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4349 = {1{`RANDOM}};
  _T_2365_re = _RAND_4349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4350 = {1{`RANDOM}};
  _T_2365_im = _RAND_4350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4351 = {1{`RANDOM}};
  _T_2366_re = _RAND_4351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4352 = {1{`RANDOM}};
  _T_2366_im = _RAND_4352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4353 = {1{`RANDOM}};
  _T_2367_re = _RAND_4353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4354 = {1{`RANDOM}};
  _T_2367_im = _RAND_4354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4355 = {1{`RANDOM}};
  _T_2368_re = _RAND_4355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4356 = {1{`RANDOM}};
  _T_2368_im = _RAND_4356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4357 = {1{`RANDOM}};
  _T_2369_re = _RAND_4357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4358 = {1{`RANDOM}};
  _T_2369_im = _RAND_4358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4359 = {1{`RANDOM}};
  _T_2370_re = _RAND_4359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4360 = {1{`RANDOM}};
  _T_2370_im = _RAND_4360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4361 = {1{`RANDOM}};
  _T_2371_re = _RAND_4361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4362 = {1{`RANDOM}};
  _T_2371_im = _RAND_4362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4363 = {1{`RANDOM}};
  _T_2372_re = _RAND_4363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4364 = {1{`RANDOM}};
  _T_2372_im = _RAND_4364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4365 = {1{`RANDOM}};
  _T_2373_re = _RAND_4365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4366 = {1{`RANDOM}};
  _T_2373_im = _RAND_4366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4367 = {1{`RANDOM}};
  _T_2374_re = _RAND_4367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4368 = {1{`RANDOM}};
  _T_2374_im = _RAND_4368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4369 = {1{`RANDOM}};
  _T_2375_re = _RAND_4369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4370 = {1{`RANDOM}};
  _T_2375_im = _RAND_4370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4371 = {1{`RANDOM}};
  _T_2376_re = _RAND_4371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4372 = {1{`RANDOM}};
  _T_2376_im = _RAND_4372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4373 = {1{`RANDOM}};
  _T_2377_re = _RAND_4373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4374 = {1{`RANDOM}};
  _T_2377_im = _RAND_4374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4375 = {1{`RANDOM}};
  _T_2378_re = _RAND_4375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4376 = {1{`RANDOM}};
  _T_2378_im = _RAND_4376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4377 = {1{`RANDOM}};
  _T_2379_re = _RAND_4377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4378 = {1{`RANDOM}};
  _T_2379_im = _RAND_4378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4379 = {1{`RANDOM}};
  _T_2380_re = _RAND_4379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4380 = {1{`RANDOM}};
  _T_2380_im = _RAND_4380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4381 = {1{`RANDOM}};
  _T_2381_re = _RAND_4381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4382 = {1{`RANDOM}};
  _T_2381_im = _RAND_4382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4383 = {1{`RANDOM}};
  _T_2382_re = _RAND_4383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4384 = {1{`RANDOM}};
  _T_2382_im = _RAND_4384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4385 = {1{`RANDOM}};
  _T_2383_re = _RAND_4385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4386 = {1{`RANDOM}};
  _T_2383_im = _RAND_4386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4387 = {1{`RANDOM}};
  _T_2384_re = _RAND_4387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4388 = {1{`RANDOM}};
  _T_2384_im = _RAND_4388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4389 = {1{`RANDOM}};
  _T_2385_re = _RAND_4389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4390 = {1{`RANDOM}};
  _T_2385_im = _RAND_4390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4391 = {1{`RANDOM}};
  _T_2386_re = _RAND_4391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4392 = {1{`RANDOM}};
  _T_2386_im = _RAND_4392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4393 = {1{`RANDOM}};
  _T_2387_re = _RAND_4393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4394 = {1{`RANDOM}};
  _T_2387_im = _RAND_4394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4395 = {1{`RANDOM}};
  _T_2388_re = _RAND_4395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4396 = {1{`RANDOM}};
  _T_2388_im = _RAND_4396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4397 = {1{`RANDOM}};
  _T_2389_re = _RAND_4397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4398 = {1{`RANDOM}};
  _T_2389_im = _RAND_4398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4399 = {1{`RANDOM}};
  _T_2390_re = _RAND_4399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4400 = {1{`RANDOM}};
  _T_2390_im = _RAND_4400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4401 = {1{`RANDOM}};
  _T_2391_re = _RAND_4401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4402 = {1{`RANDOM}};
  _T_2391_im = _RAND_4402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4403 = {1{`RANDOM}};
  _T_2392_re = _RAND_4403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4404 = {1{`RANDOM}};
  _T_2392_im = _RAND_4404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4405 = {1{`RANDOM}};
  _T_2393_re = _RAND_4405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4406 = {1{`RANDOM}};
  _T_2393_im = _RAND_4406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4407 = {1{`RANDOM}};
  _T_2394_re = _RAND_4407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4408 = {1{`RANDOM}};
  _T_2394_im = _RAND_4408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4409 = {1{`RANDOM}};
  _T_2395_re = _RAND_4409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4410 = {1{`RANDOM}};
  _T_2395_im = _RAND_4410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4411 = {1{`RANDOM}};
  _T_2396_re = _RAND_4411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4412 = {1{`RANDOM}};
  _T_2396_im = _RAND_4412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4413 = {1{`RANDOM}};
  _T_2397_re = _RAND_4413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4414 = {1{`RANDOM}};
  _T_2397_im = _RAND_4414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4415 = {1{`RANDOM}};
  _T_2398_re = _RAND_4415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4416 = {1{`RANDOM}};
  _T_2398_im = _RAND_4416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4417 = {1{`RANDOM}};
  _T_2399_re = _RAND_4417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4418 = {1{`RANDOM}};
  _T_2399_im = _RAND_4418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4419 = {1{`RANDOM}};
  _T_2400_re = _RAND_4419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4420 = {1{`RANDOM}};
  _T_2400_im = _RAND_4420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4421 = {1{`RANDOM}};
  _T_2401_re = _RAND_4421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4422 = {1{`RANDOM}};
  _T_2401_im = _RAND_4422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4423 = {1{`RANDOM}};
  _T_2402_re = _RAND_4423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4424 = {1{`RANDOM}};
  _T_2402_im = _RAND_4424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4425 = {1{`RANDOM}};
  _T_2403_re = _RAND_4425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4426 = {1{`RANDOM}};
  _T_2403_im = _RAND_4426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4427 = {1{`RANDOM}};
  _T_2404_re = _RAND_4427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4428 = {1{`RANDOM}};
  _T_2404_im = _RAND_4428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4429 = {1{`RANDOM}};
  _T_2405_re = _RAND_4429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4430 = {1{`RANDOM}};
  _T_2405_im = _RAND_4430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4431 = {1{`RANDOM}};
  _T_2406_re = _RAND_4431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4432 = {1{`RANDOM}};
  _T_2406_im = _RAND_4432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4433 = {1{`RANDOM}};
  _T_2407_re = _RAND_4433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4434 = {1{`RANDOM}};
  _T_2407_im = _RAND_4434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4435 = {1{`RANDOM}};
  _T_2408_re = _RAND_4435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4436 = {1{`RANDOM}};
  _T_2408_im = _RAND_4436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4437 = {1{`RANDOM}};
  _T_2409_re = _RAND_4437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4438 = {1{`RANDOM}};
  _T_2409_im = _RAND_4438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4439 = {1{`RANDOM}};
  _T_2410_re = _RAND_4439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4440 = {1{`RANDOM}};
  _T_2410_im = _RAND_4440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4441 = {1{`RANDOM}};
  _T_2411_re = _RAND_4441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4442 = {1{`RANDOM}};
  _T_2411_im = _RAND_4442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4443 = {1{`RANDOM}};
  _T_2412_re = _RAND_4443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4444 = {1{`RANDOM}};
  _T_2412_im = _RAND_4444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4445 = {1{`RANDOM}};
  _T_2413_re = _RAND_4445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4446 = {1{`RANDOM}};
  _T_2413_im = _RAND_4446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4447 = {1{`RANDOM}};
  _T_2414_re = _RAND_4447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4448 = {1{`RANDOM}};
  _T_2414_im = _RAND_4448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4449 = {1{`RANDOM}};
  _T_2415_re = _RAND_4449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4450 = {1{`RANDOM}};
  _T_2415_im = _RAND_4450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4451 = {1{`RANDOM}};
  _T_2416_re = _RAND_4451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4452 = {1{`RANDOM}};
  _T_2416_im = _RAND_4452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4453 = {1{`RANDOM}};
  _T_2417_re = _RAND_4453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4454 = {1{`RANDOM}};
  _T_2417_im = _RAND_4454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4455 = {1{`RANDOM}};
  _T_2418_re = _RAND_4455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4456 = {1{`RANDOM}};
  _T_2418_im = _RAND_4456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4457 = {1{`RANDOM}};
  _T_2419_re = _RAND_4457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4458 = {1{`RANDOM}};
  _T_2419_im = _RAND_4458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4459 = {1{`RANDOM}};
  _T_2420_re = _RAND_4459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4460 = {1{`RANDOM}};
  _T_2420_im = _RAND_4460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4461 = {1{`RANDOM}};
  _T_2421_re = _RAND_4461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4462 = {1{`RANDOM}};
  _T_2421_im = _RAND_4462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4463 = {1{`RANDOM}};
  _T_2422_re = _RAND_4463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4464 = {1{`RANDOM}};
  _T_2422_im = _RAND_4464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4465 = {1{`RANDOM}};
  _T_2423_re = _RAND_4465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4466 = {1{`RANDOM}};
  _T_2423_im = _RAND_4466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4467 = {1{`RANDOM}};
  _T_2424_re = _RAND_4467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4468 = {1{`RANDOM}};
  _T_2424_im = _RAND_4468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4469 = {1{`RANDOM}};
  _T_2425_re = _RAND_4469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4470 = {1{`RANDOM}};
  _T_2425_im = _RAND_4470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4471 = {1{`RANDOM}};
  _T_2426_re = _RAND_4471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4472 = {1{`RANDOM}};
  _T_2426_im = _RAND_4472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4473 = {1{`RANDOM}};
  _T_2427_re = _RAND_4473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4474 = {1{`RANDOM}};
  _T_2427_im = _RAND_4474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4475 = {1{`RANDOM}};
  _T_2428_re = _RAND_4475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4476 = {1{`RANDOM}};
  _T_2428_im = _RAND_4476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4477 = {1{`RANDOM}};
  _T_2429_re = _RAND_4477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4478 = {1{`RANDOM}};
  _T_2429_im = _RAND_4478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4479 = {1{`RANDOM}};
  _T_2430_re = _RAND_4479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4480 = {1{`RANDOM}};
  _T_2430_im = _RAND_4480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4481 = {1{`RANDOM}};
  _T_2431_re = _RAND_4481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4482 = {1{`RANDOM}};
  _T_2431_im = _RAND_4482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4483 = {1{`RANDOM}};
  _T_2432_re = _RAND_4483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4484 = {1{`RANDOM}};
  _T_2432_im = _RAND_4484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4485 = {1{`RANDOM}};
  _T_2433_re = _RAND_4485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4486 = {1{`RANDOM}};
  _T_2433_im = _RAND_4486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4487 = {1{`RANDOM}};
  _T_2434_re = _RAND_4487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4488 = {1{`RANDOM}};
  _T_2434_im = _RAND_4488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4489 = {1{`RANDOM}};
  _T_2435_re = _RAND_4489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4490 = {1{`RANDOM}};
  _T_2435_im = _RAND_4490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4491 = {1{`RANDOM}};
  _T_2436_re = _RAND_4491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4492 = {1{`RANDOM}};
  _T_2436_im = _RAND_4492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4493 = {1{`RANDOM}};
  _T_2437_re = _RAND_4493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4494 = {1{`RANDOM}};
  _T_2437_im = _RAND_4494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4495 = {1{`RANDOM}};
  _T_2438_re = _RAND_4495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4496 = {1{`RANDOM}};
  _T_2438_im = _RAND_4496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4497 = {1{`RANDOM}};
  _T_2439_re = _RAND_4497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4498 = {1{`RANDOM}};
  _T_2439_im = _RAND_4498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4499 = {1{`RANDOM}};
  _T_2440_re = _RAND_4499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4500 = {1{`RANDOM}};
  _T_2440_im = _RAND_4500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4501 = {1{`RANDOM}};
  _T_2441_re = _RAND_4501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4502 = {1{`RANDOM}};
  _T_2441_im = _RAND_4502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4503 = {1{`RANDOM}};
  _T_2442_re = _RAND_4503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4504 = {1{`RANDOM}};
  _T_2442_im = _RAND_4504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4505 = {1{`RANDOM}};
  _T_2443_re = _RAND_4505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4506 = {1{`RANDOM}};
  _T_2443_im = _RAND_4506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4507 = {1{`RANDOM}};
  _T_2444_re = _RAND_4507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4508 = {1{`RANDOM}};
  _T_2444_im = _RAND_4508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4509 = {1{`RANDOM}};
  _T_2445_re = _RAND_4509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4510 = {1{`RANDOM}};
  _T_2445_im = _RAND_4510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4511 = {1{`RANDOM}};
  _T_2446_re = _RAND_4511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4512 = {1{`RANDOM}};
  _T_2446_im = _RAND_4512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4513 = {1{`RANDOM}};
  _T_2447_re = _RAND_4513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4514 = {1{`RANDOM}};
  _T_2447_im = _RAND_4514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4515 = {1{`RANDOM}};
  _T_2448_re = _RAND_4515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4516 = {1{`RANDOM}};
  _T_2448_im = _RAND_4516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4517 = {1{`RANDOM}};
  _T_2449_re = _RAND_4517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4518 = {1{`RANDOM}};
  _T_2449_im = _RAND_4518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4519 = {1{`RANDOM}};
  _T_2450_re = _RAND_4519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4520 = {1{`RANDOM}};
  _T_2450_im = _RAND_4520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4521 = {1{`RANDOM}};
  _T_2451_re = _RAND_4521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4522 = {1{`RANDOM}};
  _T_2451_im = _RAND_4522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4523 = {1{`RANDOM}};
  _T_2452_re = _RAND_4523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4524 = {1{`RANDOM}};
  _T_2452_im = _RAND_4524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4525 = {1{`RANDOM}};
  _T_2453_re = _RAND_4525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4526 = {1{`RANDOM}};
  _T_2453_im = _RAND_4526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4527 = {1{`RANDOM}};
  _T_2454_re = _RAND_4527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4528 = {1{`RANDOM}};
  _T_2454_im = _RAND_4528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4529 = {1{`RANDOM}};
  _T_2455_re = _RAND_4529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4530 = {1{`RANDOM}};
  _T_2455_im = _RAND_4530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4531 = {1{`RANDOM}};
  _T_2456_re = _RAND_4531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4532 = {1{`RANDOM}};
  _T_2456_im = _RAND_4532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4533 = {1{`RANDOM}};
  _T_2457_re = _RAND_4533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4534 = {1{`RANDOM}};
  _T_2457_im = _RAND_4534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4535 = {1{`RANDOM}};
  _T_2458_re = _RAND_4535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4536 = {1{`RANDOM}};
  _T_2458_im = _RAND_4536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4537 = {1{`RANDOM}};
  _T_2459_re = _RAND_4537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4538 = {1{`RANDOM}};
  _T_2459_im = _RAND_4538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4539 = {1{`RANDOM}};
  _T_2460_re = _RAND_4539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4540 = {1{`RANDOM}};
  _T_2460_im = _RAND_4540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4541 = {1{`RANDOM}};
  _T_2461_re = _RAND_4541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4542 = {1{`RANDOM}};
  _T_2461_im = _RAND_4542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4543 = {1{`RANDOM}};
  _T_2462_re = _RAND_4543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4544 = {1{`RANDOM}};
  _T_2462_im = _RAND_4544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4545 = {1{`RANDOM}};
  _T_2463_re = _RAND_4545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4546 = {1{`RANDOM}};
  _T_2463_im = _RAND_4546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4547 = {1{`RANDOM}};
  _T_2464_re = _RAND_4547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4548 = {1{`RANDOM}};
  _T_2464_im = _RAND_4548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4549 = {1{`RANDOM}};
  _T_2465_re = _RAND_4549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4550 = {1{`RANDOM}};
  _T_2465_im = _RAND_4550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4551 = {1{`RANDOM}};
  _T_2466_re = _RAND_4551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4552 = {1{`RANDOM}};
  _T_2466_im = _RAND_4552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4553 = {1{`RANDOM}};
  _T_2467_re = _RAND_4553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4554 = {1{`RANDOM}};
  _T_2467_im = _RAND_4554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4555 = {1{`RANDOM}};
  _T_2468_re = _RAND_4555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4556 = {1{`RANDOM}};
  _T_2468_im = _RAND_4556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4557 = {1{`RANDOM}};
  _T_2469_re = _RAND_4557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4558 = {1{`RANDOM}};
  _T_2469_im = _RAND_4558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4559 = {1{`RANDOM}};
  _T_2470_re = _RAND_4559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4560 = {1{`RANDOM}};
  _T_2470_im = _RAND_4560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4561 = {1{`RANDOM}};
  _T_2471_re = _RAND_4561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4562 = {1{`RANDOM}};
  _T_2471_im = _RAND_4562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4563 = {1{`RANDOM}};
  _T_2472_re = _RAND_4563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4564 = {1{`RANDOM}};
  _T_2472_im = _RAND_4564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4565 = {1{`RANDOM}};
  _T_2473_re = _RAND_4565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4566 = {1{`RANDOM}};
  _T_2473_im = _RAND_4566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4567 = {1{`RANDOM}};
  _T_2474_re = _RAND_4567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4568 = {1{`RANDOM}};
  _T_2474_im = _RAND_4568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4569 = {1{`RANDOM}};
  _T_2475_re = _RAND_4569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4570 = {1{`RANDOM}};
  _T_2475_im = _RAND_4570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4571 = {1{`RANDOM}};
  _T_2476_re = _RAND_4571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4572 = {1{`RANDOM}};
  _T_2476_im = _RAND_4572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4573 = {1{`RANDOM}};
  _T_2477_re = _RAND_4573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4574 = {1{`RANDOM}};
  _T_2477_im = _RAND_4574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4575 = {1{`RANDOM}};
  _T_2478_re = _RAND_4575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4576 = {1{`RANDOM}};
  _T_2478_im = _RAND_4576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4577 = {1{`RANDOM}};
  _T_2479_re = _RAND_4577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4578 = {1{`RANDOM}};
  _T_2479_im = _RAND_4578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4579 = {1{`RANDOM}};
  _T_2480_re = _RAND_4579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4580 = {1{`RANDOM}};
  _T_2480_im = _RAND_4580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4581 = {1{`RANDOM}};
  _T_2481_re = _RAND_4581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4582 = {1{`RANDOM}};
  _T_2481_im = _RAND_4582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4583 = {1{`RANDOM}};
  _T_2482_re = _RAND_4583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4584 = {1{`RANDOM}};
  _T_2482_im = _RAND_4584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4585 = {1{`RANDOM}};
  _T_2483_re = _RAND_4585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4586 = {1{`RANDOM}};
  _T_2483_im = _RAND_4586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4587 = {1{`RANDOM}};
  _T_2484_re = _RAND_4587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4588 = {1{`RANDOM}};
  _T_2484_im = _RAND_4588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4589 = {1{`RANDOM}};
  _T_2485_re = _RAND_4589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4590 = {1{`RANDOM}};
  _T_2485_im = _RAND_4590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4591 = {1{`RANDOM}};
  _T_2486_re = _RAND_4591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4592 = {1{`RANDOM}};
  _T_2486_im = _RAND_4592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4593 = {1{`RANDOM}};
  _T_2487_re = _RAND_4593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4594 = {1{`RANDOM}};
  _T_2487_im = _RAND_4594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4595 = {1{`RANDOM}};
  _T_2488_re = _RAND_4595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4596 = {1{`RANDOM}};
  _T_2488_im = _RAND_4596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4597 = {1{`RANDOM}};
  _T_2489_re = _RAND_4597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4598 = {1{`RANDOM}};
  _T_2489_im = _RAND_4598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4599 = {1{`RANDOM}};
  _T_2490_re = _RAND_4599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4600 = {1{`RANDOM}};
  _T_2490_im = _RAND_4600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4601 = {1{`RANDOM}};
  _T_2491_re = _RAND_4601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4602 = {1{`RANDOM}};
  _T_2491_im = _RAND_4602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4603 = {1{`RANDOM}};
  _T_2492_re = _RAND_4603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4604 = {1{`RANDOM}};
  _T_2492_im = _RAND_4604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4605 = {1{`RANDOM}};
  _T_2493_re = _RAND_4605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4606 = {1{`RANDOM}};
  _T_2493_im = _RAND_4606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4607 = {1{`RANDOM}};
  _T_2494_re = _RAND_4607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4608 = {1{`RANDOM}};
  _T_2494_im = _RAND_4608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4609 = {1{`RANDOM}};
  _T_2495_re = _RAND_4609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4610 = {1{`RANDOM}};
  _T_2495_im = _RAND_4610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4611 = {1{`RANDOM}};
  _T_2496_re = _RAND_4611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4612 = {1{`RANDOM}};
  _T_2496_im = _RAND_4612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4613 = {1{`RANDOM}};
  _T_2497_re = _RAND_4613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4614 = {1{`RANDOM}};
  _T_2497_im = _RAND_4614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4615 = {1{`RANDOM}};
  _T_2507_re = _RAND_4615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4616 = {1{`RANDOM}};
  _T_2507_im = _RAND_4616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4617 = {1{`RANDOM}};
  _T_2508_re = _RAND_4617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4618 = {1{`RANDOM}};
  _T_2508_im = _RAND_4618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4619 = {1{`RANDOM}};
  _T_2509_re = _RAND_4619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4620 = {1{`RANDOM}};
  _T_2509_im = _RAND_4620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4621 = {1{`RANDOM}};
  _T_2510_re = _RAND_4621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4622 = {1{`RANDOM}};
  _T_2510_im = _RAND_4622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4623 = {1{`RANDOM}};
  _T_2511_re = _RAND_4623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4624 = {1{`RANDOM}};
  _T_2511_im = _RAND_4624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4625 = {1{`RANDOM}};
  _T_2512_re = _RAND_4625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4626 = {1{`RANDOM}};
  _T_2512_im = _RAND_4626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4627 = {1{`RANDOM}};
  _T_2513_re = _RAND_4627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4628 = {1{`RANDOM}};
  _T_2513_im = _RAND_4628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4629 = {1{`RANDOM}};
  _T_2514_re = _RAND_4629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4630 = {1{`RANDOM}};
  _T_2514_im = _RAND_4630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4631 = {1{`RANDOM}};
  _T_2515_re = _RAND_4631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4632 = {1{`RANDOM}};
  _T_2515_im = _RAND_4632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4633 = {1{`RANDOM}};
  _T_2516_re = _RAND_4633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4634 = {1{`RANDOM}};
  _T_2516_im = _RAND_4634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4635 = {1{`RANDOM}};
  _T_2517_re = _RAND_4635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4636 = {1{`RANDOM}};
  _T_2517_im = _RAND_4636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4637 = {1{`RANDOM}};
  _T_2518_re = _RAND_4637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4638 = {1{`RANDOM}};
  _T_2518_im = _RAND_4638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4639 = {1{`RANDOM}};
  _T_2519_re = _RAND_4639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4640 = {1{`RANDOM}};
  _T_2519_im = _RAND_4640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4641 = {1{`RANDOM}};
  _T_2520_re = _RAND_4641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4642 = {1{`RANDOM}};
  _T_2520_im = _RAND_4642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4643 = {1{`RANDOM}};
  _T_2521_re = _RAND_4643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4644 = {1{`RANDOM}};
  _T_2521_im = _RAND_4644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4645 = {1{`RANDOM}};
  _T_2522_re = _RAND_4645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4646 = {1{`RANDOM}};
  _T_2522_im = _RAND_4646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4647 = {1{`RANDOM}};
  _T_2523_re = _RAND_4647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4648 = {1{`RANDOM}};
  _T_2523_im = _RAND_4648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4649 = {1{`RANDOM}};
  _T_2524_re = _RAND_4649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4650 = {1{`RANDOM}};
  _T_2524_im = _RAND_4650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4651 = {1{`RANDOM}};
  _T_2525_re = _RAND_4651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4652 = {1{`RANDOM}};
  _T_2525_im = _RAND_4652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4653 = {1{`RANDOM}};
  _T_2526_re = _RAND_4653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4654 = {1{`RANDOM}};
  _T_2526_im = _RAND_4654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4655 = {1{`RANDOM}};
  _T_2527_re = _RAND_4655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4656 = {1{`RANDOM}};
  _T_2527_im = _RAND_4656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4657 = {1{`RANDOM}};
  _T_2528_re = _RAND_4657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4658 = {1{`RANDOM}};
  _T_2528_im = _RAND_4658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4659 = {1{`RANDOM}};
  _T_2529_re = _RAND_4659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4660 = {1{`RANDOM}};
  _T_2529_im = _RAND_4660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4661 = {1{`RANDOM}};
  _T_2530_re = _RAND_4661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4662 = {1{`RANDOM}};
  _T_2530_im = _RAND_4662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4663 = {1{`RANDOM}};
  _T_2531_re = _RAND_4663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4664 = {1{`RANDOM}};
  _T_2531_im = _RAND_4664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4665 = {1{`RANDOM}};
  _T_2532_re = _RAND_4665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4666 = {1{`RANDOM}};
  _T_2532_im = _RAND_4666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4667 = {1{`RANDOM}};
  _T_2533_re = _RAND_4667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4668 = {1{`RANDOM}};
  _T_2533_im = _RAND_4668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4669 = {1{`RANDOM}};
  _T_2534_re = _RAND_4669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4670 = {1{`RANDOM}};
  _T_2534_im = _RAND_4670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4671 = {1{`RANDOM}};
  _T_2535_re = _RAND_4671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4672 = {1{`RANDOM}};
  _T_2535_im = _RAND_4672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4673 = {1{`RANDOM}};
  _T_2536_re = _RAND_4673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4674 = {1{`RANDOM}};
  _T_2536_im = _RAND_4674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4675 = {1{`RANDOM}};
  _T_2537_re = _RAND_4675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4676 = {1{`RANDOM}};
  _T_2537_im = _RAND_4676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4677 = {1{`RANDOM}};
  _T_2538_re = _RAND_4677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4678 = {1{`RANDOM}};
  _T_2538_im = _RAND_4678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4679 = {1{`RANDOM}};
  _T_2539_re = _RAND_4679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4680 = {1{`RANDOM}};
  _T_2539_im = _RAND_4680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4681 = {1{`RANDOM}};
  _T_2540_re = _RAND_4681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4682 = {1{`RANDOM}};
  _T_2540_im = _RAND_4682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4683 = {1{`RANDOM}};
  _T_2541_re = _RAND_4683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4684 = {1{`RANDOM}};
  _T_2541_im = _RAND_4684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4685 = {1{`RANDOM}};
  _T_2542_re = _RAND_4685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4686 = {1{`RANDOM}};
  _T_2542_im = _RAND_4686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4687 = {1{`RANDOM}};
  _T_2543_re = _RAND_4687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4688 = {1{`RANDOM}};
  _T_2543_im = _RAND_4688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4689 = {1{`RANDOM}};
  _T_2544_re = _RAND_4689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4690 = {1{`RANDOM}};
  _T_2544_im = _RAND_4690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4691 = {1{`RANDOM}};
  _T_2545_re = _RAND_4691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4692 = {1{`RANDOM}};
  _T_2545_im = _RAND_4692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4693 = {1{`RANDOM}};
  _T_2546_re = _RAND_4693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4694 = {1{`RANDOM}};
  _T_2546_im = _RAND_4694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4695 = {1{`RANDOM}};
  _T_2547_re = _RAND_4695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4696 = {1{`RANDOM}};
  _T_2547_im = _RAND_4696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4697 = {1{`RANDOM}};
  _T_2548_re = _RAND_4697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4698 = {1{`RANDOM}};
  _T_2548_im = _RAND_4698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4699 = {1{`RANDOM}};
  _T_2549_re = _RAND_4699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4700 = {1{`RANDOM}};
  _T_2549_im = _RAND_4700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4701 = {1{`RANDOM}};
  _T_2550_re = _RAND_4701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4702 = {1{`RANDOM}};
  _T_2550_im = _RAND_4702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4703 = {1{`RANDOM}};
  _T_2551_re = _RAND_4703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4704 = {1{`RANDOM}};
  _T_2551_im = _RAND_4704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4705 = {1{`RANDOM}};
  _T_2552_re = _RAND_4705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4706 = {1{`RANDOM}};
  _T_2552_im = _RAND_4706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4707 = {1{`RANDOM}};
  _T_2553_re = _RAND_4707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4708 = {1{`RANDOM}};
  _T_2553_im = _RAND_4708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4709 = {1{`RANDOM}};
  _T_2554_re = _RAND_4709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4710 = {1{`RANDOM}};
  _T_2554_im = _RAND_4710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4711 = {1{`RANDOM}};
  _T_2555_re = _RAND_4711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4712 = {1{`RANDOM}};
  _T_2555_im = _RAND_4712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4713 = {1{`RANDOM}};
  _T_2556_re = _RAND_4713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4714 = {1{`RANDOM}};
  _T_2556_im = _RAND_4714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4715 = {1{`RANDOM}};
  _T_2557_re = _RAND_4715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4716 = {1{`RANDOM}};
  _T_2557_im = _RAND_4716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4717 = {1{`RANDOM}};
  _T_2558_re = _RAND_4717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4718 = {1{`RANDOM}};
  _T_2558_im = _RAND_4718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4719 = {1{`RANDOM}};
  _T_2559_re = _RAND_4719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4720 = {1{`RANDOM}};
  _T_2559_im = _RAND_4720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4721 = {1{`RANDOM}};
  _T_2560_re = _RAND_4721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4722 = {1{`RANDOM}};
  _T_2560_im = _RAND_4722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4723 = {1{`RANDOM}};
  _T_2561_re = _RAND_4723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4724 = {1{`RANDOM}};
  _T_2561_im = _RAND_4724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4725 = {1{`RANDOM}};
  _T_2562_re = _RAND_4725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4726 = {1{`RANDOM}};
  _T_2562_im = _RAND_4726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4727 = {1{`RANDOM}};
  _T_2563_re = _RAND_4727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4728 = {1{`RANDOM}};
  _T_2563_im = _RAND_4728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4729 = {1{`RANDOM}};
  _T_2564_re = _RAND_4729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4730 = {1{`RANDOM}};
  _T_2564_im = _RAND_4730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4731 = {1{`RANDOM}};
  _T_2565_re = _RAND_4731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4732 = {1{`RANDOM}};
  _T_2565_im = _RAND_4732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4733 = {1{`RANDOM}};
  _T_2566_re = _RAND_4733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4734 = {1{`RANDOM}};
  _T_2566_im = _RAND_4734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4735 = {1{`RANDOM}};
  _T_2567_re = _RAND_4735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4736 = {1{`RANDOM}};
  _T_2567_im = _RAND_4736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4737 = {1{`RANDOM}};
  _T_2568_re = _RAND_4737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4738 = {1{`RANDOM}};
  _T_2568_im = _RAND_4738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4739 = {1{`RANDOM}};
  _T_2569_re = _RAND_4739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4740 = {1{`RANDOM}};
  _T_2569_im = _RAND_4740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4741 = {1{`RANDOM}};
  _T_2570_re = _RAND_4741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4742 = {1{`RANDOM}};
  _T_2570_im = _RAND_4742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4743 = {1{`RANDOM}};
  _T_2571_re = _RAND_4743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4744 = {1{`RANDOM}};
  _T_2571_im = _RAND_4744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4745 = {1{`RANDOM}};
  _T_2572_re = _RAND_4745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4746 = {1{`RANDOM}};
  _T_2572_im = _RAND_4746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4747 = {1{`RANDOM}};
  _T_2573_re = _RAND_4747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4748 = {1{`RANDOM}};
  _T_2573_im = _RAND_4748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4749 = {1{`RANDOM}};
  _T_2574_re = _RAND_4749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4750 = {1{`RANDOM}};
  _T_2574_im = _RAND_4750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4751 = {1{`RANDOM}};
  _T_2575_re = _RAND_4751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4752 = {1{`RANDOM}};
  _T_2575_im = _RAND_4752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4753 = {1{`RANDOM}};
  _T_2576_re = _RAND_4753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4754 = {1{`RANDOM}};
  _T_2576_im = _RAND_4754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4755 = {1{`RANDOM}};
  _T_2577_re = _RAND_4755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4756 = {1{`RANDOM}};
  _T_2577_im = _RAND_4756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4757 = {1{`RANDOM}};
  _T_2578_re = _RAND_4757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4758 = {1{`RANDOM}};
  _T_2578_im = _RAND_4758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4759 = {1{`RANDOM}};
  _T_2579_re = _RAND_4759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4760 = {1{`RANDOM}};
  _T_2579_im = _RAND_4760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4761 = {1{`RANDOM}};
  _T_2580_re = _RAND_4761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4762 = {1{`RANDOM}};
  _T_2580_im = _RAND_4762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4763 = {1{`RANDOM}};
  _T_2581_re = _RAND_4763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4764 = {1{`RANDOM}};
  _T_2581_im = _RAND_4764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4765 = {1{`RANDOM}};
  _T_2582_re = _RAND_4765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4766 = {1{`RANDOM}};
  _T_2582_im = _RAND_4766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4767 = {1{`RANDOM}};
  _T_2583_re = _RAND_4767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4768 = {1{`RANDOM}};
  _T_2583_im = _RAND_4768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4769 = {1{`RANDOM}};
  _T_2584_re = _RAND_4769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4770 = {1{`RANDOM}};
  _T_2584_im = _RAND_4770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4771 = {1{`RANDOM}};
  _T_2585_re = _RAND_4771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4772 = {1{`RANDOM}};
  _T_2585_im = _RAND_4772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4773 = {1{`RANDOM}};
  _T_2586_re = _RAND_4773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4774 = {1{`RANDOM}};
  _T_2586_im = _RAND_4774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4775 = {1{`RANDOM}};
  _T_2587_re = _RAND_4775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4776 = {1{`RANDOM}};
  _T_2587_im = _RAND_4776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4777 = {1{`RANDOM}};
  _T_2588_re = _RAND_4777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4778 = {1{`RANDOM}};
  _T_2588_im = _RAND_4778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4779 = {1{`RANDOM}};
  _T_2589_re = _RAND_4779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4780 = {1{`RANDOM}};
  _T_2589_im = _RAND_4780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4781 = {1{`RANDOM}};
  _T_2590_re = _RAND_4781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4782 = {1{`RANDOM}};
  _T_2590_im = _RAND_4782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4783 = {1{`RANDOM}};
  _T_2591_re = _RAND_4783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4784 = {1{`RANDOM}};
  _T_2591_im = _RAND_4784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4785 = {1{`RANDOM}};
  _T_2592_re = _RAND_4785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4786 = {1{`RANDOM}};
  _T_2592_im = _RAND_4786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4787 = {1{`RANDOM}};
  _T_2593_re = _RAND_4787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4788 = {1{`RANDOM}};
  _T_2593_im = _RAND_4788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4789 = {1{`RANDOM}};
  _T_2594_re = _RAND_4789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4790 = {1{`RANDOM}};
  _T_2594_im = _RAND_4790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4791 = {1{`RANDOM}};
  _T_2595_re = _RAND_4791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4792 = {1{`RANDOM}};
  _T_2595_im = _RAND_4792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4793 = {1{`RANDOM}};
  _T_2596_re = _RAND_4793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4794 = {1{`RANDOM}};
  _T_2596_im = _RAND_4794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4795 = {1{`RANDOM}};
  _T_2597_re = _RAND_4795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4796 = {1{`RANDOM}};
  _T_2597_im = _RAND_4796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4797 = {1{`RANDOM}};
  _T_2598_re = _RAND_4797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4798 = {1{`RANDOM}};
  _T_2598_im = _RAND_4798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4799 = {1{`RANDOM}};
  _T_2599_re = _RAND_4799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4800 = {1{`RANDOM}};
  _T_2599_im = _RAND_4800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4801 = {1{`RANDOM}};
  _T_2600_re = _RAND_4801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4802 = {1{`RANDOM}};
  _T_2600_im = _RAND_4802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4803 = {1{`RANDOM}};
  _T_2601_re = _RAND_4803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4804 = {1{`RANDOM}};
  _T_2601_im = _RAND_4804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4805 = {1{`RANDOM}};
  _T_2602_re = _RAND_4805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4806 = {1{`RANDOM}};
  _T_2602_im = _RAND_4806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4807 = {1{`RANDOM}};
  _T_2603_re = _RAND_4807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4808 = {1{`RANDOM}};
  _T_2603_im = _RAND_4808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4809 = {1{`RANDOM}};
  _T_2604_re = _RAND_4809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4810 = {1{`RANDOM}};
  _T_2604_im = _RAND_4810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4811 = {1{`RANDOM}};
  _T_2605_re = _RAND_4811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4812 = {1{`RANDOM}};
  _T_2605_im = _RAND_4812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4813 = {1{`RANDOM}};
  _T_2606_re = _RAND_4813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4814 = {1{`RANDOM}};
  _T_2606_im = _RAND_4814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4815 = {1{`RANDOM}};
  _T_2607_re = _RAND_4815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4816 = {1{`RANDOM}};
  _T_2607_im = _RAND_4816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4817 = {1{`RANDOM}};
  _T_2608_re = _RAND_4817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4818 = {1{`RANDOM}};
  _T_2608_im = _RAND_4818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4819 = {1{`RANDOM}};
  _T_2609_re = _RAND_4819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4820 = {1{`RANDOM}};
  _T_2609_im = _RAND_4820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4821 = {1{`RANDOM}};
  _T_2610_re = _RAND_4821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4822 = {1{`RANDOM}};
  _T_2610_im = _RAND_4822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4823 = {1{`RANDOM}};
  _T_2611_re = _RAND_4823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4824 = {1{`RANDOM}};
  _T_2611_im = _RAND_4824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4825 = {1{`RANDOM}};
  _T_2612_re = _RAND_4825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4826 = {1{`RANDOM}};
  _T_2612_im = _RAND_4826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4827 = {1{`RANDOM}};
  _T_2613_re = _RAND_4827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4828 = {1{`RANDOM}};
  _T_2613_im = _RAND_4828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4829 = {1{`RANDOM}};
  _T_2614_re = _RAND_4829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4830 = {1{`RANDOM}};
  _T_2614_im = _RAND_4830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4831 = {1{`RANDOM}};
  _T_2615_re = _RAND_4831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4832 = {1{`RANDOM}};
  _T_2615_im = _RAND_4832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4833 = {1{`RANDOM}};
  _T_2616_re = _RAND_4833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4834 = {1{`RANDOM}};
  _T_2616_im = _RAND_4834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4835 = {1{`RANDOM}};
  _T_2617_re = _RAND_4835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4836 = {1{`RANDOM}};
  _T_2617_im = _RAND_4836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4837 = {1{`RANDOM}};
  _T_2618_re = _RAND_4837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4838 = {1{`RANDOM}};
  _T_2618_im = _RAND_4838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4839 = {1{`RANDOM}};
  _T_2619_re = _RAND_4839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4840 = {1{`RANDOM}};
  _T_2619_im = _RAND_4840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4841 = {1{`RANDOM}};
  _T_2620_re = _RAND_4841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4842 = {1{`RANDOM}};
  _T_2620_im = _RAND_4842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4843 = {1{`RANDOM}};
  _T_2621_re = _RAND_4843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4844 = {1{`RANDOM}};
  _T_2621_im = _RAND_4844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4845 = {1{`RANDOM}};
  _T_2622_re = _RAND_4845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4846 = {1{`RANDOM}};
  _T_2622_im = _RAND_4846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4847 = {1{`RANDOM}};
  _T_2623_re = _RAND_4847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4848 = {1{`RANDOM}};
  _T_2623_im = _RAND_4848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4849 = {1{`RANDOM}};
  _T_2624_re = _RAND_4849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4850 = {1{`RANDOM}};
  _T_2624_im = _RAND_4850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4851 = {1{`RANDOM}};
  _T_2625_re = _RAND_4851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4852 = {1{`RANDOM}};
  _T_2625_im = _RAND_4852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4853 = {1{`RANDOM}};
  _T_2626_re = _RAND_4853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4854 = {1{`RANDOM}};
  _T_2626_im = _RAND_4854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4855 = {1{`RANDOM}};
  _T_2627_re = _RAND_4855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4856 = {1{`RANDOM}};
  _T_2627_im = _RAND_4856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4857 = {1{`RANDOM}};
  _T_2628_re = _RAND_4857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4858 = {1{`RANDOM}};
  _T_2628_im = _RAND_4858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4859 = {1{`RANDOM}};
  _T_2629_re = _RAND_4859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4860 = {1{`RANDOM}};
  _T_2629_im = _RAND_4860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4861 = {1{`RANDOM}};
  _T_2630_re = _RAND_4861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4862 = {1{`RANDOM}};
  _T_2630_im = _RAND_4862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4863 = {1{`RANDOM}};
  _T_2631_re = _RAND_4863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4864 = {1{`RANDOM}};
  _T_2631_im = _RAND_4864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4865 = {1{`RANDOM}};
  _T_2632_re = _RAND_4865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4866 = {1{`RANDOM}};
  _T_2632_im = _RAND_4866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4867 = {1{`RANDOM}};
  _T_2633_re = _RAND_4867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4868 = {1{`RANDOM}};
  _T_2633_im = _RAND_4868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4869 = {1{`RANDOM}};
  _T_2634_re = _RAND_4869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4870 = {1{`RANDOM}};
  _T_2634_im = _RAND_4870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4871 = {1{`RANDOM}};
  _T_2635_re = _RAND_4871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4872 = {1{`RANDOM}};
  _T_2635_im = _RAND_4872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4873 = {1{`RANDOM}};
  _T_2636_re = _RAND_4873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4874 = {1{`RANDOM}};
  _T_2636_im = _RAND_4874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4875 = {1{`RANDOM}};
  _T_2637_re = _RAND_4875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4876 = {1{`RANDOM}};
  _T_2637_im = _RAND_4876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4877 = {1{`RANDOM}};
  _T_2638_re = _RAND_4877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4878 = {1{`RANDOM}};
  _T_2638_im = _RAND_4878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4879 = {1{`RANDOM}};
  _T_2639_re = _RAND_4879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4880 = {1{`RANDOM}};
  _T_2639_im = _RAND_4880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4881 = {1{`RANDOM}};
  _T_2640_re = _RAND_4881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4882 = {1{`RANDOM}};
  _T_2640_im = _RAND_4882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4883 = {1{`RANDOM}};
  _T_2641_re = _RAND_4883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4884 = {1{`RANDOM}};
  _T_2641_im = _RAND_4884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4885 = {1{`RANDOM}};
  _T_2642_re = _RAND_4885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4886 = {1{`RANDOM}};
  _T_2642_im = _RAND_4886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4887 = {1{`RANDOM}};
  _T_2643_re = _RAND_4887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4888 = {1{`RANDOM}};
  _T_2643_im = _RAND_4888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4889 = {1{`RANDOM}};
  _T_2644_re = _RAND_4889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4890 = {1{`RANDOM}};
  _T_2644_im = _RAND_4890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4891 = {1{`RANDOM}};
  _T_2645_re = _RAND_4891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4892 = {1{`RANDOM}};
  _T_2645_im = _RAND_4892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4893 = {1{`RANDOM}};
  _T_2646_re = _RAND_4893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4894 = {1{`RANDOM}};
  _T_2646_im = _RAND_4894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4895 = {1{`RANDOM}};
  _T_2647_re = _RAND_4895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4896 = {1{`RANDOM}};
  _T_2647_im = _RAND_4896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4897 = {1{`RANDOM}};
  _T_2648_re = _RAND_4897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4898 = {1{`RANDOM}};
  _T_2648_im = _RAND_4898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4899 = {1{`RANDOM}};
  _T_2649_re = _RAND_4899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4900 = {1{`RANDOM}};
  _T_2649_im = _RAND_4900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4901 = {1{`RANDOM}};
  _T_2650_re = _RAND_4901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4902 = {1{`RANDOM}};
  _T_2650_im = _RAND_4902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4903 = {1{`RANDOM}};
  _T_2651_re = _RAND_4903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4904 = {1{`RANDOM}};
  _T_2651_im = _RAND_4904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4905 = {1{`RANDOM}};
  _T_2652_re = _RAND_4905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4906 = {1{`RANDOM}};
  _T_2652_im = _RAND_4906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4907 = {1{`RANDOM}};
  _T_2653_re = _RAND_4907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4908 = {1{`RANDOM}};
  _T_2653_im = _RAND_4908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4909 = {1{`RANDOM}};
  _T_2654_re = _RAND_4909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4910 = {1{`RANDOM}};
  _T_2654_im = _RAND_4910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4911 = {1{`RANDOM}};
  _T_2655_re = _RAND_4911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4912 = {1{`RANDOM}};
  _T_2655_im = _RAND_4912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4913 = {1{`RANDOM}};
  _T_2656_re = _RAND_4913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4914 = {1{`RANDOM}};
  _T_2656_im = _RAND_4914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4915 = {1{`RANDOM}};
  _T_2657_re = _RAND_4915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4916 = {1{`RANDOM}};
  _T_2657_im = _RAND_4916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4917 = {1{`RANDOM}};
  _T_2658_re = _RAND_4917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4918 = {1{`RANDOM}};
  _T_2658_im = _RAND_4918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4919 = {1{`RANDOM}};
  _T_2659_re = _RAND_4919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4920 = {1{`RANDOM}};
  _T_2659_im = _RAND_4920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4921 = {1{`RANDOM}};
  _T_2660_re = _RAND_4921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4922 = {1{`RANDOM}};
  _T_2660_im = _RAND_4922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4923 = {1{`RANDOM}};
  _T_2661_re = _RAND_4923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4924 = {1{`RANDOM}};
  _T_2661_im = _RAND_4924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4925 = {1{`RANDOM}};
  _T_2662_re = _RAND_4925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4926 = {1{`RANDOM}};
  _T_2662_im = _RAND_4926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4927 = {1{`RANDOM}};
  _T_2663_re = _RAND_4927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4928 = {1{`RANDOM}};
  _T_2663_im = _RAND_4928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4929 = {1{`RANDOM}};
  _T_2664_re = _RAND_4929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4930 = {1{`RANDOM}};
  _T_2664_im = _RAND_4930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4931 = {1{`RANDOM}};
  _T_2665_re = _RAND_4931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4932 = {1{`RANDOM}};
  _T_2665_im = _RAND_4932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4933 = {1{`RANDOM}};
  _T_2666_re = _RAND_4933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4934 = {1{`RANDOM}};
  _T_2666_im = _RAND_4934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4935 = {1{`RANDOM}};
  _T_2667_re = _RAND_4935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4936 = {1{`RANDOM}};
  _T_2667_im = _RAND_4936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4937 = {1{`RANDOM}};
  _T_2668_re = _RAND_4937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4938 = {1{`RANDOM}};
  _T_2668_im = _RAND_4938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4939 = {1{`RANDOM}};
  _T_2669_re = _RAND_4939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4940 = {1{`RANDOM}};
  _T_2669_im = _RAND_4940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4941 = {1{`RANDOM}};
  _T_2670_re = _RAND_4941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4942 = {1{`RANDOM}};
  _T_2670_im = _RAND_4942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4943 = {1{`RANDOM}};
  _T_2671_re = _RAND_4943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4944 = {1{`RANDOM}};
  _T_2671_im = _RAND_4944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4945 = {1{`RANDOM}};
  _T_2672_re = _RAND_4945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4946 = {1{`RANDOM}};
  _T_2672_im = _RAND_4946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4947 = {1{`RANDOM}};
  _T_2673_re = _RAND_4947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4948 = {1{`RANDOM}};
  _T_2673_im = _RAND_4948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4949 = {1{`RANDOM}};
  _T_2674_re = _RAND_4949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4950 = {1{`RANDOM}};
  _T_2674_im = _RAND_4950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4951 = {1{`RANDOM}};
  _T_2675_re = _RAND_4951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4952 = {1{`RANDOM}};
  _T_2675_im = _RAND_4952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4953 = {1{`RANDOM}};
  _T_2676_re = _RAND_4953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4954 = {1{`RANDOM}};
  _T_2676_im = _RAND_4954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4955 = {1{`RANDOM}};
  _T_2677_re = _RAND_4955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4956 = {1{`RANDOM}};
  _T_2677_im = _RAND_4956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4957 = {1{`RANDOM}};
  _T_2678_re = _RAND_4957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4958 = {1{`RANDOM}};
  _T_2678_im = _RAND_4958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4959 = {1{`RANDOM}};
  _T_2679_re = _RAND_4959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4960 = {1{`RANDOM}};
  _T_2679_im = _RAND_4960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4961 = {1{`RANDOM}};
  _T_2680_re = _RAND_4961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4962 = {1{`RANDOM}};
  _T_2680_im = _RAND_4962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4963 = {1{`RANDOM}};
  _T_2681_re = _RAND_4963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4964 = {1{`RANDOM}};
  _T_2681_im = _RAND_4964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4965 = {1{`RANDOM}};
  _T_2682_re = _RAND_4965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4966 = {1{`RANDOM}};
  _T_2682_im = _RAND_4966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4967 = {1{`RANDOM}};
  _T_2683_re = _RAND_4967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4968 = {1{`RANDOM}};
  _T_2683_im = _RAND_4968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4969 = {1{`RANDOM}};
  _T_2684_re = _RAND_4969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4970 = {1{`RANDOM}};
  _T_2684_im = _RAND_4970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4971 = {1{`RANDOM}};
  _T_2685_re = _RAND_4971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4972 = {1{`RANDOM}};
  _T_2685_im = _RAND_4972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4973 = {1{`RANDOM}};
  _T_2686_re = _RAND_4973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4974 = {1{`RANDOM}};
  _T_2686_im = _RAND_4974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4975 = {1{`RANDOM}};
  _T_2687_re = _RAND_4975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4976 = {1{`RANDOM}};
  _T_2687_im = _RAND_4976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4977 = {1{`RANDOM}};
  _T_2688_re = _RAND_4977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4978 = {1{`RANDOM}};
  _T_2688_im = _RAND_4978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4979 = {1{`RANDOM}};
  _T_2689_re = _RAND_4979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4980 = {1{`RANDOM}};
  _T_2689_im = _RAND_4980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4981 = {1{`RANDOM}};
  _T_2690_re = _RAND_4981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4982 = {1{`RANDOM}};
  _T_2690_im = _RAND_4982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4983 = {1{`RANDOM}};
  _T_2691_re = _RAND_4983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4984 = {1{`RANDOM}};
  _T_2691_im = _RAND_4984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4985 = {1{`RANDOM}};
  _T_2692_re = _RAND_4985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4986 = {1{`RANDOM}};
  _T_2692_im = _RAND_4986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4987 = {1{`RANDOM}};
  _T_2693_re = _RAND_4987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4988 = {1{`RANDOM}};
  _T_2693_im = _RAND_4988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4989 = {1{`RANDOM}};
  _T_2694_re = _RAND_4989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4990 = {1{`RANDOM}};
  _T_2694_im = _RAND_4990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4991 = {1{`RANDOM}};
  _T_2695_re = _RAND_4991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4992 = {1{`RANDOM}};
  _T_2695_im = _RAND_4992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4993 = {1{`RANDOM}};
  _T_2696_re = _RAND_4993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4994 = {1{`RANDOM}};
  _T_2696_im = _RAND_4994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4995 = {1{`RANDOM}};
  _T_2697_re = _RAND_4995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4996 = {1{`RANDOM}};
  _T_2697_im = _RAND_4996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4997 = {1{`RANDOM}};
  _T_2698_re = _RAND_4997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4998 = {1{`RANDOM}};
  _T_2698_im = _RAND_4998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4999 = {1{`RANDOM}};
  _T_2699_re = _RAND_4999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5000 = {1{`RANDOM}};
  _T_2699_im = _RAND_5000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5001 = {1{`RANDOM}};
  _T_2700_re = _RAND_5001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5002 = {1{`RANDOM}};
  _T_2700_im = _RAND_5002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5003 = {1{`RANDOM}};
  _T_2701_re = _RAND_5003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5004 = {1{`RANDOM}};
  _T_2701_im = _RAND_5004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5005 = {1{`RANDOM}};
  _T_2702_re = _RAND_5005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5006 = {1{`RANDOM}};
  _T_2702_im = _RAND_5006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5007 = {1{`RANDOM}};
  _T_2703_re = _RAND_5007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5008 = {1{`RANDOM}};
  _T_2703_im = _RAND_5008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5009 = {1{`RANDOM}};
  _T_2704_re = _RAND_5009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5010 = {1{`RANDOM}};
  _T_2704_im = _RAND_5010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5011 = {1{`RANDOM}};
  _T_2705_re = _RAND_5011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5012 = {1{`RANDOM}};
  _T_2705_im = _RAND_5012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5013 = {1{`RANDOM}};
  _T_2706_re = _RAND_5013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5014 = {1{`RANDOM}};
  _T_2706_im = _RAND_5014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5015 = {1{`RANDOM}};
  _T_2707_re = _RAND_5015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5016 = {1{`RANDOM}};
  _T_2707_im = _RAND_5016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5017 = {1{`RANDOM}};
  _T_2708_re = _RAND_5017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5018 = {1{`RANDOM}};
  _T_2708_im = _RAND_5018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5019 = {1{`RANDOM}};
  _T_2709_re = _RAND_5019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5020 = {1{`RANDOM}};
  _T_2709_im = _RAND_5020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5021 = {1{`RANDOM}};
  _T_2710_re = _RAND_5021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5022 = {1{`RANDOM}};
  _T_2710_im = _RAND_5022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5023 = {1{`RANDOM}};
  _T_2711_re = _RAND_5023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5024 = {1{`RANDOM}};
  _T_2711_im = _RAND_5024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5025 = {1{`RANDOM}};
  _T_2712_re = _RAND_5025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5026 = {1{`RANDOM}};
  _T_2712_im = _RAND_5026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5027 = {1{`RANDOM}};
  _T_2713_re = _RAND_5027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5028 = {1{`RANDOM}};
  _T_2713_im = _RAND_5028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5029 = {1{`RANDOM}};
  _T_2714_re = _RAND_5029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5030 = {1{`RANDOM}};
  _T_2714_im = _RAND_5030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5031 = {1{`RANDOM}};
  _T_2715_re = _RAND_5031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5032 = {1{`RANDOM}};
  _T_2715_im = _RAND_5032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5033 = {1{`RANDOM}};
  _T_2716_re = _RAND_5033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5034 = {1{`RANDOM}};
  _T_2716_im = _RAND_5034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5035 = {1{`RANDOM}};
  _T_2717_re = _RAND_5035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5036 = {1{`RANDOM}};
  _T_2717_im = _RAND_5036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5037 = {1{`RANDOM}};
  _T_2718_re = _RAND_5037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5038 = {1{`RANDOM}};
  _T_2718_im = _RAND_5038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5039 = {1{`RANDOM}};
  _T_2719_re = _RAND_5039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5040 = {1{`RANDOM}};
  _T_2719_im = _RAND_5040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5041 = {1{`RANDOM}};
  _T_2720_re = _RAND_5041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5042 = {1{`RANDOM}};
  _T_2720_im = _RAND_5042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5043 = {1{`RANDOM}};
  _T_2721_re = _RAND_5043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5044 = {1{`RANDOM}};
  _T_2721_im = _RAND_5044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5045 = {1{`RANDOM}};
  _T_2722_re = _RAND_5045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5046 = {1{`RANDOM}};
  _T_2722_im = _RAND_5046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5047 = {1{`RANDOM}};
  _T_2723_re = _RAND_5047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5048 = {1{`RANDOM}};
  _T_2723_im = _RAND_5048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5049 = {1{`RANDOM}};
  _T_2724_re = _RAND_5049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5050 = {1{`RANDOM}};
  _T_2724_im = _RAND_5050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5051 = {1{`RANDOM}};
  _T_2725_re = _RAND_5051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5052 = {1{`RANDOM}};
  _T_2725_im = _RAND_5052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5053 = {1{`RANDOM}};
  _T_2726_re = _RAND_5053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5054 = {1{`RANDOM}};
  _T_2726_im = _RAND_5054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5055 = {1{`RANDOM}};
  _T_2727_re = _RAND_5055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5056 = {1{`RANDOM}};
  _T_2727_im = _RAND_5056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5057 = {1{`RANDOM}};
  _T_2728_re = _RAND_5057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5058 = {1{`RANDOM}};
  _T_2728_im = _RAND_5058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5059 = {1{`RANDOM}};
  _T_2729_re = _RAND_5059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5060 = {1{`RANDOM}};
  _T_2729_im = _RAND_5060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5061 = {1{`RANDOM}};
  _T_2730_re = _RAND_5061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5062 = {1{`RANDOM}};
  _T_2730_im = _RAND_5062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5063 = {1{`RANDOM}};
  _T_2731_re = _RAND_5063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5064 = {1{`RANDOM}};
  _T_2731_im = _RAND_5064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5065 = {1{`RANDOM}};
  _T_2732_re = _RAND_5065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5066 = {1{`RANDOM}};
  _T_2732_im = _RAND_5066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5067 = {1{`RANDOM}};
  _T_2733_re = _RAND_5067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5068 = {1{`RANDOM}};
  _T_2733_im = _RAND_5068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5069 = {1{`RANDOM}};
  _T_2734_re = _RAND_5069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5070 = {1{`RANDOM}};
  _T_2734_im = _RAND_5070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5071 = {1{`RANDOM}};
  _T_2735_re = _RAND_5071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5072 = {1{`RANDOM}};
  _T_2735_im = _RAND_5072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5073 = {1{`RANDOM}};
  _T_2736_re = _RAND_5073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5074 = {1{`RANDOM}};
  _T_2736_im = _RAND_5074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5075 = {1{`RANDOM}};
  _T_2737_re = _RAND_5075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5076 = {1{`RANDOM}};
  _T_2737_im = _RAND_5076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5077 = {1{`RANDOM}};
  _T_2738_re = _RAND_5077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5078 = {1{`RANDOM}};
  _T_2738_im = _RAND_5078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5079 = {1{`RANDOM}};
  _T_2739_re = _RAND_5079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5080 = {1{`RANDOM}};
  _T_2739_im = _RAND_5080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5081 = {1{`RANDOM}};
  _T_2740_re = _RAND_5081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5082 = {1{`RANDOM}};
  _T_2740_im = _RAND_5082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5083 = {1{`RANDOM}};
  _T_2741_re = _RAND_5083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5084 = {1{`RANDOM}};
  _T_2741_im = _RAND_5084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5085 = {1{`RANDOM}};
  _T_2742_re = _RAND_5085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5086 = {1{`RANDOM}};
  _T_2742_im = _RAND_5086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5087 = {1{`RANDOM}};
  _T_2743_re = _RAND_5087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5088 = {1{`RANDOM}};
  _T_2743_im = _RAND_5088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5089 = {1{`RANDOM}};
  _T_2744_re = _RAND_5089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5090 = {1{`RANDOM}};
  _T_2744_im = _RAND_5090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5091 = {1{`RANDOM}};
  _T_2745_re = _RAND_5091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5092 = {1{`RANDOM}};
  _T_2745_im = _RAND_5092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5093 = {1{`RANDOM}};
  _T_2746_re = _RAND_5093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5094 = {1{`RANDOM}};
  _T_2746_im = _RAND_5094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5095 = {1{`RANDOM}};
  _T_2747_re = _RAND_5095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5096 = {1{`RANDOM}};
  _T_2747_im = _RAND_5096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5097 = {1{`RANDOM}};
  _T_2748_re = _RAND_5097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5098 = {1{`RANDOM}};
  _T_2748_im = _RAND_5098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5099 = {1{`RANDOM}};
  _T_2749_re = _RAND_5099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5100 = {1{`RANDOM}};
  _T_2749_im = _RAND_5100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5101 = {1{`RANDOM}};
  _T_2750_re = _RAND_5101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5102 = {1{`RANDOM}};
  _T_2750_im = _RAND_5102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5103 = {1{`RANDOM}};
  _T_2751_re = _RAND_5103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5104 = {1{`RANDOM}};
  _T_2751_im = _RAND_5104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5105 = {1{`RANDOM}};
  _T_2752_re = _RAND_5105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5106 = {1{`RANDOM}};
  _T_2752_im = _RAND_5106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5107 = {1{`RANDOM}};
  _T_2753_re = _RAND_5107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5108 = {1{`RANDOM}};
  _T_2753_im = _RAND_5108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5109 = {1{`RANDOM}};
  _T_2754_re = _RAND_5109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5110 = {1{`RANDOM}};
  _T_2754_im = _RAND_5110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5111 = {1{`RANDOM}};
  _T_2755_re = _RAND_5111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5112 = {1{`RANDOM}};
  _T_2755_im = _RAND_5112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5113 = {1{`RANDOM}};
  _T_2756_re = _RAND_5113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5114 = {1{`RANDOM}};
  _T_2756_im = _RAND_5114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5115 = {1{`RANDOM}};
  _T_2757_re = _RAND_5115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5116 = {1{`RANDOM}};
  _T_2757_im = _RAND_5116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5117 = {1{`RANDOM}};
  _T_2758_re = _RAND_5117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5118 = {1{`RANDOM}};
  _T_2758_im = _RAND_5118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5119 = {1{`RANDOM}};
  _T_2759_re = _RAND_5119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5120 = {1{`RANDOM}};
  _T_2759_im = _RAND_5120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5121 = {1{`RANDOM}};
  _T_2760_re = _RAND_5121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5122 = {1{`RANDOM}};
  _T_2760_im = _RAND_5122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5123 = {1{`RANDOM}};
  _T_2761_re = _RAND_5123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5124 = {1{`RANDOM}};
  _T_2761_im = _RAND_5124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5125 = {1{`RANDOM}};
  _T_2762_re = _RAND_5125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5126 = {1{`RANDOM}};
  _T_2762_im = _RAND_5126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5127 = {1{`RANDOM}};
  _T_2765_re = _RAND_5127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5128 = {1{`RANDOM}};
  _T_2765_im = _RAND_5128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5129 = {1{`RANDOM}};
  _T_2766_re = _RAND_5129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5130 = {1{`RANDOM}};
  _T_2766_im = _RAND_5130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5131 = {1{`RANDOM}};
  _T_2767_re = _RAND_5131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5132 = {1{`RANDOM}};
  _T_2767_im = _RAND_5132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5133 = {1{`RANDOM}};
  _T_2768_re = _RAND_5133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5134 = {1{`RANDOM}};
  _T_2768_im = _RAND_5134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5135 = {1{`RANDOM}};
  _T_2769_re = _RAND_5135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5136 = {1{`RANDOM}};
  _T_2769_im = _RAND_5136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5137 = {1{`RANDOM}};
  _T_2770_re = _RAND_5137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5138 = {1{`RANDOM}};
  _T_2770_im = _RAND_5138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5139 = {1{`RANDOM}};
  _T_2771_re = _RAND_5139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5140 = {1{`RANDOM}};
  _T_2771_im = _RAND_5140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5141 = {1{`RANDOM}};
  _T_2772_re = _RAND_5141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5142 = {1{`RANDOM}};
  _T_2772_im = _RAND_5142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5143 = {1{`RANDOM}};
  _T_2773_re = _RAND_5143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5144 = {1{`RANDOM}};
  _T_2773_im = _RAND_5144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5145 = {1{`RANDOM}};
  _T_2774_re = _RAND_5145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5146 = {1{`RANDOM}};
  _T_2774_im = _RAND_5146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5147 = {1{`RANDOM}};
  _T_2775_re = _RAND_5147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5148 = {1{`RANDOM}};
  _T_2775_im = _RAND_5148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5149 = {1{`RANDOM}};
  _T_2776_re = _RAND_5149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5150 = {1{`RANDOM}};
  _T_2776_im = _RAND_5150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5151 = {1{`RANDOM}};
  _T_2777_re = _RAND_5151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5152 = {1{`RANDOM}};
  _T_2777_im = _RAND_5152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5153 = {1{`RANDOM}};
  _T_2778_re = _RAND_5153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5154 = {1{`RANDOM}};
  _T_2778_im = _RAND_5154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5155 = {1{`RANDOM}};
  _T_2779_re = _RAND_5155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5156 = {1{`RANDOM}};
  _T_2779_im = _RAND_5156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5157 = {1{`RANDOM}};
  _T_2780_re = _RAND_5157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5158 = {1{`RANDOM}};
  _T_2780_im = _RAND_5158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5159 = {1{`RANDOM}};
  _T_2781_re = _RAND_5159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5160 = {1{`RANDOM}};
  _T_2781_im = _RAND_5160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5161 = {1{`RANDOM}};
  _T_2782_re = _RAND_5161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5162 = {1{`RANDOM}};
  _T_2782_im = _RAND_5162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5163 = {1{`RANDOM}};
  _T_2783_re = _RAND_5163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5164 = {1{`RANDOM}};
  _T_2783_im = _RAND_5164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5165 = {1{`RANDOM}};
  _T_2784_re = _RAND_5165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5166 = {1{`RANDOM}};
  _T_2784_im = _RAND_5166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5167 = {1{`RANDOM}};
  _T_2785_re = _RAND_5167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5168 = {1{`RANDOM}};
  _T_2785_im = _RAND_5168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5169 = {1{`RANDOM}};
  _T_2786_re = _RAND_5169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5170 = {1{`RANDOM}};
  _T_2786_im = _RAND_5170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5171 = {1{`RANDOM}};
  _T_2787_re = _RAND_5171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5172 = {1{`RANDOM}};
  _T_2787_im = _RAND_5172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5173 = {1{`RANDOM}};
  _T_2788_re = _RAND_5173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5174 = {1{`RANDOM}};
  _T_2788_im = _RAND_5174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5175 = {1{`RANDOM}};
  _T_2789_re = _RAND_5175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5176 = {1{`RANDOM}};
  _T_2789_im = _RAND_5176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5177 = {1{`RANDOM}};
  _T_2790_re = _RAND_5177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5178 = {1{`RANDOM}};
  _T_2790_im = _RAND_5178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5179 = {1{`RANDOM}};
  _T_2791_re = _RAND_5179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5180 = {1{`RANDOM}};
  _T_2791_im = _RAND_5180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5181 = {1{`RANDOM}};
  _T_2792_re = _RAND_5181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5182 = {1{`RANDOM}};
  _T_2792_im = _RAND_5182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5183 = {1{`RANDOM}};
  _T_2793_re = _RAND_5183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5184 = {1{`RANDOM}};
  _T_2793_im = _RAND_5184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5185 = {1{`RANDOM}};
  _T_2794_re = _RAND_5185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5186 = {1{`RANDOM}};
  _T_2794_im = _RAND_5186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5187 = {1{`RANDOM}};
  _T_2795_re = _RAND_5187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5188 = {1{`RANDOM}};
  _T_2795_im = _RAND_5188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5189 = {1{`RANDOM}};
  _T_2796_re = _RAND_5189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5190 = {1{`RANDOM}};
  _T_2796_im = _RAND_5190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5191 = {1{`RANDOM}};
  _T_2797_re = _RAND_5191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5192 = {1{`RANDOM}};
  _T_2797_im = _RAND_5192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5193 = {1{`RANDOM}};
  _T_2798_re = _RAND_5193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5194 = {1{`RANDOM}};
  _T_2798_im = _RAND_5194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5195 = {1{`RANDOM}};
  _T_2799_re = _RAND_5195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5196 = {1{`RANDOM}};
  _T_2799_im = _RAND_5196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5197 = {1{`RANDOM}};
  _T_2800_re = _RAND_5197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5198 = {1{`RANDOM}};
  _T_2800_im = _RAND_5198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5199 = {1{`RANDOM}};
  _T_2801_re = _RAND_5199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5200 = {1{`RANDOM}};
  _T_2801_im = _RAND_5200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5201 = {1{`RANDOM}};
  _T_2802_re = _RAND_5201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5202 = {1{`RANDOM}};
  _T_2802_im = _RAND_5202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5203 = {1{`RANDOM}};
  _T_2803_re = _RAND_5203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5204 = {1{`RANDOM}};
  _T_2803_im = _RAND_5204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5205 = {1{`RANDOM}};
  _T_2804_re = _RAND_5205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5206 = {1{`RANDOM}};
  _T_2804_im = _RAND_5206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5207 = {1{`RANDOM}};
  _T_2805_re = _RAND_5207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5208 = {1{`RANDOM}};
  _T_2805_im = _RAND_5208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5209 = {1{`RANDOM}};
  _T_2806_re = _RAND_5209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5210 = {1{`RANDOM}};
  _T_2806_im = _RAND_5210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5211 = {1{`RANDOM}};
  _T_2807_re = _RAND_5211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5212 = {1{`RANDOM}};
  _T_2807_im = _RAND_5212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5213 = {1{`RANDOM}};
  _T_2808_re = _RAND_5213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5214 = {1{`RANDOM}};
  _T_2808_im = _RAND_5214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5215 = {1{`RANDOM}};
  _T_2809_re = _RAND_5215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5216 = {1{`RANDOM}};
  _T_2809_im = _RAND_5216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5217 = {1{`RANDOM}};
  _T_2810_re = _RAND_5217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5218 = {1{`RANDOM}};
  _T_2810_im = _RAND_5218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5219 = {1{`RANDOM}};
  _T_2811_re = _RAND_5219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5220 = {1{`RANDOM}};
  _T_2811_im = _RAND_5220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5221 = {1{`RANDOM}};
  _T_2812_re = _RAND_5221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5222 = {1{`RANDOM}};
  _T_2812_im = _RAND_5222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5223 = {1{`RANDOM}};
  _T_2813_re = _RAND_5223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5224 = {1{`RANDOM}};
  _T_2813_im = _RAND_5224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5225 = {1{`RANDOM}};
  _T_2814_re = _RAND_5225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5226 = {1{`RANDOM}};
  _T_2814_im = _RAND_5226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5227 = {1{`RANDOM}};
  _T_2815_re = _RAND_5227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5228 = {1{`RANDOM}};
  _T_2815_im = _RAND_5228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5229 = {1{`RANDOM}};
  _T_2816_re = _RAND_5229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5230 = {1{`RANDOM}};
  _T_2816_im = _RAND_5230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5231 = {1{`RANDOM}};
  _T_2817_re = _RAND_5231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5232 = {1{`RANDOM}};
  _T_2817_im = _RAND_5232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5233 = {1{`RANDOM}};
  _T_2818_re = _RAND_5233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5234 = {1{`RANDOM}};
  _T_2818_im = _RAND_5234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5235 = {1{`RANDOM}};
  _T_2819_re = _RAND_5235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5236 = {1{`RANDOM}};
  _T_2819_im = _RAND_5236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5237 = {1{`RANDOM}};
  _T_2820_re = _RAND_5237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5238 = {1{`RANDOM}};
  _T_2820_im = _RAND_5238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5239 = {1{`RANDOM}};
  _T_2821_re = _RAND_5239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5240 = {1{`RANDOM}};
  _T_2821_im = _RAND_5240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5241 = {1{`RANDOM}};
  _T_2822_re = _RAND_5241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5242 = {1{`RANDOM}};
  _T_2822_im = _RAND_5242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5243 = {1{`RANDOM}};
  _T_2823_re = _RAND_5243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5244 = {1{`RANDOM}};
  _T_2823_im = _RAND_5244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5245 = {1{`RANDOM}};
  _T_2824_re = _RAND_5245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5246 = {1{`RANDOM}};
  _T_2824_im = _RAND_5246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5247 = {1{`RANDOM}};
  _T_2825_re = _RAND_5247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5248 = {1{`RANDOM}};
  _T_2825_im = _RAND_5248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5249 = {1{`RANDOM}};
  _T_2826_re = _RAND_5249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5250 = {1{`RANDOM}};
  _T_2826_im = _RAND_5250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5251 = {1{`RANDOM}};
  _T_2827_re = _RAND_5251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5252 = {1{`RANDOM}};
  _T_2827_im = _RAND_5252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5253 = {1{`RANDOM}};
  _T_2828_re = _RAND_5253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5254 = {1{`RANDOM}};
  _T_2828_im = _RAND_5254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5255 = {1{`RANDOM}};
  _T_2829_re = _RAND_5255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5256 = {1{`RANDOM}};
  _T_2829_im = _RAND_5256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5257 = {1{`RANDOM}};
  _T_2830_re = _RAND_5257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5258 = {1{`RANDOM}};
  _T_2830_im = _RAND_5258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5259 = {1{`RANDOM}};
  _T_2831_re = _RAND_5259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5260 = {1{`RANDOM}};
  _T_2831_im = _RAND_5260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5261 = {1{`RANDOM}};
  _T_2832_re = _RAND_5261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5262 = {1{`RANDOM}};
  _T_2832_im = _RAND_5262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5263 = {1{`RANDOM}};
  _T_2833_re = _RAND_5263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5264 = {1{`RANDOM}};
  _T_2833_im = _RAND_5264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5265 = {1{`RANDOM}};
  _T_2834_re = _RAND_5265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5266 = {1{`RANDOM}};
  _T_2834_im = _RAND_5266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5267 = {1{`RANDOM}};
  _T_2835_re = _RAND_5267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5268 = {1{`RANDOM}};
  _T_2835_im = _RAND_5268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5269 = {1{`RANDOM}};
  _T_2836_re = _RAND_5269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5270 = {1{`RANDOM}};
  _T_2836_im = _RAND_5270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5271 = {1{`RANDOM}};
  _T_2837_re = _RAND_5271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5272 = {1{`RANDOM}};
  _T_2837_im = _RAND_5272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5273 = {1{`RANDOM}};
  _T_2838_re = _RAND_5273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5274 = {1{`RANDOM}};
  _T_2838_im = _RAND_5274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5275 = {1{`RANDOM}};
  _T_2839_re = _RAND_5275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5276 = {1{`RANDOM}};
  _T_2839_im = _RAND_5276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5277 = {1{`RANDOM}};
  _T_2840_re = _RAND_5277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5278 = {1{`RANDOM}};
  _T_2840_im = _RAND_5278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5279 = {1{`RANDOM}};
  _T_2841_re = _RAND_5279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5280 = {1{`RANDOM}};
  _T_2841_im = _RAND_5280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5281 = {1{`RANDOM}};
  _T_2842_re = _RAND_5281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5282 = {1{`RANDOM}};
  _T_2842_im = _RAND_5282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5283 = {1{`RANDOM}};
  _T_2843_re = _RAND_5283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5284 = {1{`RANDOM}};
  _T_2843_im = _RAND_5284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5285 = {1{`RANDOM}};
  _T_2844_re = _RAND_5285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5286 = {1{`RANDOM}};
  _T_2844_im = _RAND_5286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5287 = {1{`RANDOM}};
  _T_2845_re = _RAND_5287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5288 = {1{`RANDOM}};
  _T_2845_im = _RAND_5288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5289 = {1{`RANDOM}};
  _T_2846_re = _RAND_5289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5290 = {1{`RANDOM}};
  _T_2846_im = _RAND_5290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5291 = {1{`RANDOM}};
  _T_2847_re = _RAND_5291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5292 = {1{`RANDOM}};
  _T_2847_im = _RAND_5292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5293 = {1{`RANDOM}};
  _T_2848_re = _RAND_5293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5294 = {1{`RANDOM}};
  _T_2848_im = _RAND_5294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5295 = {1{`RANDOM}};
  _T_2849_re = _RAND_5295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5296 = {1{`RANDOM}};
  _T_2849_im = _RAND_5296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5297 = {1{`RANDOM}};
  _T_2850_re = _RAND_5297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5298 = {1{`RANDOM}};
  _T_2850_im = _RAND_5298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5299 = {1{`RANDOM}};
  _T_2851_re = _RAND_5299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5300 = {1{`RANDOM}};
  _T_2851_im = _RAND_5300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5301 = {1{`RANDOM}};
  _T_2852_re = _RAND_5301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5302 = {1{`RANDOM}};
  _T_2852_im = _RAND_5302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5303 = {1{`RANDOM}};
  _T_2853_re = _RAND_5303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5304 = {1{`RANDOM}};
  _T_2853_im = _RAND_5304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5305 = {1{`RANDOM}};
  _T_2854_re = _RAND_5305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5306 = {1{`RANDOM}};
  _T_2854_im = _RAND_5306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5307 = {1{`RANDOM}};
  _T_2855_re = _RAND_5307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5308 = {1{`RANDOM}};
  _T_2855_im = _RAND_5308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5309 = {1{`RANDOM}};
  _T_2856_re = _RAND_5309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5310 = {1{`RANDOM}};
  _T_2856_im = _RAND_5310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5311 = {1{`RANDOM}};
  _T_2857_re = _RAND_5311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5312 = {1{`RANDOM}};
  _T_2857_im = _RAND_5312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5313 = {1{`RANDOM}};
  _T_2858_re = _RAND_5313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5314 = {1{`RANDOM}};
  _T_2858_im = _RAND_5314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5315 = {1{`RANDOM}};
  _T_2859_re = _RAND_5315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5316 = {1{`RANDOM}};
  _T_2859_im = _RAND_5316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5317 = {1{`RANDOM}};
  _T_2860_re = _RAND_5317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5318 = {1{`RANDOM}};
  _T_2860_im = _RAND_5318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5319 = {1{`RANDOM}};
  _T_2861_re = _RAND_5319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5320 = {1{`RANDOM}};
  _T_2861_im = _RAND_5320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5321 = {1{`RANDOM}};
  _T_2862_re = _RAND_5321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5322 = {1{`RANDOM}};
  _T_2862_im = _RAND_5322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5323 = {1{`RANDOM}};
  _T_2863_re = _RAND_5323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5324 = {1{`RANDOM}};
  _T_2863_im = _RAND_5324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5325 = {1{`RANDOM}};
  _T_2864_re = _RAND_5325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5326 = {1{`RANDOM}};
  _T_2864_im = _RAND_5326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5327 = {1{`RANDOM}};
  _T_2865_re = _RAND_5327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5328 = {1{`RANDOM}};
  _T_2865_im = _RAND_5328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5329 = {1{`RANDOM}};
  _T_2866_re = _RAND_5329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5330 = {1{`RANDOM}};
  _T_2866_im = _RAND_5330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5331 = {1{`RANDOM}};
  _T_2867_re = _RAND_5331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5332 = {1{`RANDOM}};
  _T_2867_im = _RAND_5332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5333 = {1{`RANDOM}};
  _T_2868_re = _RAND_5333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5334 = {1{`RANDOM}};
  _T_2868_im = _RAND_5334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5335 = {1{`RANDOM}};
  _T_2869_re = _RAND_5335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5336 = {1{`RANDOM}};
  _T_2869_im = _RAND_5336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5337 = {1{`RANDOM}};
  _T_2870_re = _RAND_5337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5338 = {1{`RANDOM}};
  _T_2870_im = _RAND_5338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5339 = {1{`RANDOM}};
  _T_2871_re = _RAND_5339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5340 = {1{`RANDOM}};
  _T_2871_im = _RAND_5340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5341 = {1{`RANDOM}};
  _T_2872_re = _RAND_5341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5342 = {1{`RANDOM}};
  _T_2872_im = _RAND_5342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5343 = {1{`RANDOM}};
  _T_2873_re = _RAND_5343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5344 = {1{`RANDOM}};
  _T_2873_im = _RAND_5344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5345 = {1{`RANDOM}};
  _T_2874_re = _RAND_5345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5346 = {1{`RANDOM}};
  _T_2874_im = _RAND_5346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5347 = {1{`RANDOM}};
  _T_2875_re = _RAND_5347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5348 = {1{`RANDOM}};
  _T_2875_im = _RAND_5348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5349 = {1{`RANDOM}};
  _T_2876_re = _RAND_5349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5350 = {1{`RANDOM}};
  _T_2876_im = _RAND_5350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5351 = {1{`RANDOM}};
  _T_2877_re = _RAND_5351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5352 = {1{`RANDOM}};
  _T_2877_im = _RAND_5352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5353 = {1{`RANDOM}};
  _T_2878_re = _RAND_5353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5354 = {1{`RANDOM}};
  _T_2878_im = _RAND_5354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5355 = {1{`RANDOM}};
  _T_2879_re = _RAND_5355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5356 = {1{`RANDOM}};
  _T_2879_im = _RAND_5356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5357 = {1{`RANDOM}};
  _T_2880_re = _RAND_5357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5358 = {1{`RANDOM}};
  _T_2880_im = _RAND_5358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5359 = {1{`RANDOM}};
  _T_2881_re = _RAND_5359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5360 = {1{`RANDOM}};
  _T_2881_im = _RAND_5360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5361 = {1{`RANDOM}};
  _T_2882_re = _RAND_5361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5362 = {1{`RANDOM}};
  _T_2882_im = _RAND_5362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5363 = {1{`RANDOM}};
  _T_2883_re = _RAND_5363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5364 = {1{`RANDOM}};
  _T_2883_im = _RAND_5364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5365 = {1{`RANDOM}};
  _T_2884_re = _RAND_5365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5366 = {1{`RANDOM}};
  _T_2884_im = _RAND_5366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5367 = {1{`RANDOM}};
  _T_2885_re = _RAND_5367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5368 = {1{`RANDOM}};
  _T_2885_im = _RAND_5368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5369 = {1{`RANDOM}};
  _T_2886_re = _RAND_5369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5370 = {1{`RANDOM}};
  _T_2886_im = _RAND_5370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5371 = {1{`RANDOM}};
  _T_2887_re = _RAND_5371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5372 = {1{`RANDOM}};
  _T_2887_im = _RAND_5372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5373 = {1{`RANDOM}};
  _T_2888_re = _RAND_5373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5374 = {1{`RANDOM}};
  _T_2888_im = _RAND_5374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5375 = {1{`RANDOM}};
  _T_2889_re = _RAND_5375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5376 = {1{`RANDOM}};
  _T_2889_im = _RAND_5376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5377 = {1{`RANDOM}};
  _T_2890_re = _RAND_5377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5378 = {1{`RANDOM}};
  _T_2890_im = _RAND_5378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5379 = {1{`RANDOM}};
  _T_2891_re = _RAND_5379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5380 = {1{`RANDOM}};
  _T_2891_im = _RAND_5380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5381 = {1{`RANDOM}};
  _T_2892_re = _RAND_5381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5382 = {1{`RANDOM}};
  _T_2892_im = _RAND_5382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5383 = {1{`RANDOM}};
  _T_2902_re = _RAND_5383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5384 = {1{`RANDOM}};
  _T_2902_im = _RAND_5384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5385 = {1{`RANDOM}};
  _T_2903_re = _RAND_5385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5386 = {1{`RANDOM}};
  _T_2903_im = _RAND_5386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5387 = {1{`RANDOM}};
  _T_2904_re = _RAND_5387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5388 = {1{`RANDOM}};
  _T_2904_im = _RAND_5388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5389 = {1{`RANDOM}};
  _T_2905_re = _RAND_5389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5390 = {1{`RANDOM}};
  _T_2905_im = _RAND_5390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5391 = {1{`RANDOM}};
  _T_2906_re = _RAND_5391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5392 = {1{`RANDOM}};
  _T_2906_im = _RAND_5392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5393 = {1{`RANDOM}};
  _T_2907_re = _RAND_5393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5394 = {1{`RANDOM}};
  _T_2907_im = _RAND_5394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5395 = {1{`RANDOM}};
  _T_2908_re = _RAND_5395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5396 = {1{`RANDOM}};
  _T_2908_im = _RAND_5396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5397 = {1{`RANDOM}};
  _T_2909_re = _RAND_5397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5398 = {1{`RANDOM}};
  _T_2909_im = _RAND_5398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5399 = {1{`RANDOM}};
  _T_2910_re = _RAND_5399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5400 = {1{`RANDOM}};
  _T_2910_im = _RAND_5400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5401 = {1{`RANDOM}};
  _T_2911_re = _RAND_5401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5402 = {1{`RANDOM}};
  _T_2911_im = _RAND_5402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5403 = {1{`RANDOM}};
  _T_2912_re = _RAND_5403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5404 = {1{`RANDOM}};
  _T_2912_im = _RAND_5404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5405 = {1{`RANDOM}};
  _T_2913_re = _RAND_5405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5406 = {1{`RANDOM}};
  _T_2913_im = _RAND_5406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5407 = {1{`RANDOM}};
  _T_2914_re = _RAND_5407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5408 = {1{`RANDOM}};
  _T_2914_im = _RAND_5408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5409 = {1{`RANDOM}};
  _T_2915_re = _RAND_5409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5410 = {1{`RANDOM}};
  _T_2915_im = _RAND_5410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5411 = {1{`RANDOM}};
  _T_2916_re = _RAND_5411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5412 = {1{`RANDOM}};
  _T_2916_im = _RAND_5412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5413 = {1{`RANDOM}};
  _T_2917_re = _RAND_5413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5414 = {1{`RANDOM}};
  _T_2917_im = _RAND_5414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5415 = {1{`RANDOM}};
  _T_2918_re = _RAND_5415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5416 = {1{`RANDOM}};
  _T_2918_im = _RAND_5416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5417 = {1{`RANDOM}};
  _T_2919_re = _RAND_5417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5418 = {1{`RANDOM}};
  _T_2919_im = _RAND_5418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5419 = {1{`RANDOM}};
  _T_2920_re = _RAND_5419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5420 = {1{`RANDOM}};
  _T_2920_im = _RAND_5420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5421 = {1{`RANDOM}};
  _T_2921_re = _RAND_5421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5422 = {1{`RANDOM}};
  _T_2921_im = _RAND_5422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5423 = {1{`RANDOM}};
  _T_2922_re = _RAND_5423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5424 = {1{`RANDOM}};
  _T_2922_im = _RAND_5424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5425 = {1{`RANDOM}};
  _T_2923_re = _RAND_5425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5426 = {1{`RANDOM}};
  _T_2923_im = _RAND_5426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5427 = {1{`RANDOM}};
  _T_2924_re = _RAND_5427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5428 = {1{`RANDOM}};
  _T_2924_im = _RAND_5428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5429 = {1{`RANDOM}};
  _T_2925_re = _RAND_5429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5430 = {1{`RANDOM}};
  _T_2925_im = _RAND_5430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5431 = {1{`RANDOM}};
  _T_2926_re = _RAND_5431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5432 = {1{`RANDOM}};
  _T_2926_im = _RAND_5432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5433 = {1{`RANDOM}};
  _T_2927_re = _RAND_5433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5434 = {1{`RANDOM}};
  _T_2927_im = _RAND_5434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5435 = {1{`RANDOM}};
  _T_2928_re = _RAND_5435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5436 = {1{`RANDOM}};
  _T_2928_im = _RAND_5436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5437 = {1{`RANDOM}};
  _T_2929_re = _RAND_5437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5438 = {1{`RANDOM}};
  _T_2929_im = _RAND_5438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5439 = {1{`RANDOM}};
  _T_2930_re = _RAND_5439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5440 = {1{`RANDOM}};
  _T_2930_im = _RAND_5440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5441 = {1{`RANDOM}};
  _T_2931_re = _RAND_5441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5442 = {1{`RANDOM}};
  _T_2931_im = _RAND_5442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5443 = {1{`RANDOM}};
  _T_2932_re = _RAND_5443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5444 = {1{`RANDOM}};
  _T_2932_im = _RAND_5444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5445 = {1{`RANDOM}};
  _T_2933_re = _RAND_5445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5446 = {1{`RANDOM}};
  _T_2933_im = _RAND_5446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5447 = {1{`RANDOM}};
  _T_2934_re = _RAND_5447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5448 = {1{`RANDOM}};
  _T_2934_im = _RAND_5448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5449 = {1{`RANDOM}};
  _T_2935_re = _RAND_5449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5450 = {1{`RANDOM}};
  _T_2935_im = _RAND_5450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5451 = {1{`RANDOM}};
  _T_2936_re = _RAND_5451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5452 = {1{`RANDOM}};
  _T_2936_im = _RAND_5452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5453 = {1{`RANDOM}};
  _T_2937_re = _RAND_5453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5454 = {1{`RANDOM}};
  _T_2937_im = _RAND_5454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5455 = {1{`RANDOM}};
  _T_2938_re = _RAND_5455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5456 = {1{`RANDOM}};
  _T_2938_im = _RAND_5456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5457 = {1{`RANDOM}};
  _T_2939_re = _RAND_5457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5458 = {1{`RANDOM}};
  _T_2939_im = _RAND_5458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5459 = {1{`RANDOM}};
  _T_2940_re = _RAND_5459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5460 = {1{`RANDOM}};
  _T_2940_im = _RAND_5460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5461 = {1{`RANDOM}};
  _T_2941_re = _RAND_5461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5462 = {1{`RANDOM}};
  _T_2941_im = _RAND_5462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5463 = {1{`RANDOM}};
  _T_2942_re = _RAND_5463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5464 = {1{`RANDOM}};
  _T_2942_im = _RAND_5464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5465 = {1{`RANDOM}};
  _T_2943_re = _RAND_5465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5466 = {1{`RANDOM}};
  _T_2943_im = _RAND_5466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5467 = {1{`RANDOM}};
  _T_2944_re = _RAND_5467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5468 = {1{`RANDOM}};
  _T_2944_im = _RAND_5468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5469 = {1{`RANDOM}};
  _T_2945_re = _RAND_5469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5470 = {1{`RANDOM}};
  _T_2945_im = _RAND_5470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5471 = {1{`RANDOM}};
  _T_2946_re = _RAND_5471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5472 = {1{`RANDOM}};
  _T_2946_im = _RAND_5472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5473 = {1{`RANDOM}};
  _T_2947_re = _RAND_5473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5474 = {1{`RANDOM}};
  _T_2947_im = _RAND_5474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5475 = {1{`RANDOM}};
  _T_2948_re = _RAND_5475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5476 = {1{`RANDOM}};
  _T_2948_im = _RAND_5476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5477 = {1{`RANDOM}};
  _T_2949_re = _RAND_5477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5478 = {1{`RANDOM}};
  _T_2949_im = _RAND_5478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5479 = {1{`RANDOM}};
  _T_2950_re = _RAND_5479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5480 = {1{`RANDOM}};
  _T_2950_im = _RAND_5480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5481 = {1{`RANDOM}};
  _T_2951_re = _RAND_5481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5482 = {1{`RANDOM}};
  _T_2951_im = _RAND_5482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5483 = {1{`RANDOM}};
  _T_2952_re = _RAND_5483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5484 = {1{`RANDOM}};
  _T_2952_im = _RAND_5484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5485 = {1{`RANDOM}};
  _T_2953_re = _RAND_5485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5486 = {1{`RANDOM}};
  _T_2953_im = _RAND_5486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5487 = {1{`RANDOM}};
  _T_2954_re = _RAND_5487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5488 = {1{`RANDOM}};
  _T_2954_im = _RAND_5488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5489 = {1{`RANDOM}};
  _T_2955_re = _RAND_5489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5490 = {1{`RANDOM}};
  _T_2955_im = _RAND_5490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5491 = {1{`RANDOM}};
  _T_2956_re = _RAND_5491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5492 = {1{`RANDOM}};
  _T_2956_im = _RAND_5492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5493 = {1{`RANDOM}};
  _T_2957_re = _RAND_5493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5494 = {1{`RANDOM}};
  _T_2957_im = _RAND_5494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5495 = {1{`RANDOM}};
  _T_2958_re = _RAND_5495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5496 = {1{`RANDOM}};
  _T_2958_im = _RAND_5496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5497 = {1{`RANDOM}};
  _T_2959_re = _RAND_5497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5498 = {1{`RANDOM}};
  _T_2959_im = _RAND_5498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5499 = {1{`RANDOM}};
  _T_2960_re = _RAND_5499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5500 = {1{`RANDOM}};
  _T_2960_im = _RAND_5500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5501 = {1{`RANDOM}};
  _T_2961_re = _RAND_5501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5502 = {1{`RANDOM}};
  _T_2961_im = _RAND_5502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5503 = {1{`RANDOM}};
  _T_2962_re = _RAND_5503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5504 = {1{`RANDOM}};
  _T_2962_im = _RAND_5504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5505 = {1{`RANDOM}};
  _T_2963_re = _RAND_5505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5506 = {1{`RANDOM}};
  _T_2963_im = _RAND_5506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5507 = {1{`RANDOM}};
  _T_2964_re = _RAND_5507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5508 = {1{`RANDOM}};
  _T_2964_im = _RAND_5508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5509 = {1{`RANDOM}};
  _T_2965_re = _RAND_5509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5510 = {1{`RANDOM}};
  _T_2965_im = _RAND_5510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5511 = {1{`RANDOM}};
  _T_2966_re = _RAND_5511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5512 = {1{`RANDOM}};
  _T_2966_im = _RAND_5512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5513 = {1{`RANDOM}};
  _T_2967_re = _RAND_5513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5514 = {1{`RANDOM}};
  _T_2967_im = _RAND_5514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5515 = {1{`RANDOM}};
  _T_2968_re = _RAND_5515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5516 = {1{`RANDOM}};
  _T_2968_im = _RAND_5516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5517 = {1{`RANDOM}};
  _T_2969_re = _RAND_5517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5518 = {1{`RANDOM}};
  _T_2969_im = _RAND_5518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5519 = {1{`RANDOM}};
  _T_2970_re = _RAND_5519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5520 = {1{`RANDOM}};
  _T_2970_im = _RAND_5520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5521 = {1{`RANDOM}};
  _T_2971_re = _RAND_5521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5522 = {1{`RANDOM}};
  _T_2971_im = _RAND_5522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5523 = {1{`RANDOM}};
  _T_2972_re = _RAND_5523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5524 = {1{`RANDOM}};
  _T_2972_im = _RAND_5524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5525 = {1{`RANDOM}};
  _T_2973_re = _RAND_5525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5526 = {1{`RANDOM}};
  _T_2973_im = _RAND_5526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5527 = {1{`RANDOM}};
  _T_2974_re = _RAND_5527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5528 = {1{`RANDOM}};
  _T_2974_im = _RAND_5528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5529 = {1{`RANDOM}};
  _T_2975_re = _RAND_5529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5530 = {1{`RANDOM}};
  _T_2975_im = _RAND_5530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5531 = {1{`RANDOM}};
  _T_2976_re = _RAND_5531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5532 = {1{`RANDOM}};
  _T_2976_im = _RAND_5532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5533 = {1{`RANDOM}};
  _T_2977_re = _RAND_5533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5534 = {1{`RANDOM}};
  _T_2977_im = _RAND_5534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5535 = {1{`RANDOM}};
  _T_2978_re = _RAND_5535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5536 = {1{`RANDOM}};
  _T_2978_im = _RAND_5536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5537 = {1{`RANDOM}};
  _T_2979_re = _RAND_5537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5538 = {1{`RANDOM}};
  _T_2979_im = _RAND_5538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5539 = {1{`RANDOM}};
  _T_2980_re = _RAND_5539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5540 = {1{`RANDOM}};
  _T_2980_im = _RAND_5540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5541 = {1{`RANDOM}};
  _T_2981_re = _RAND_5541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5542 = {1{`RANDOM}};
  _T_2981_im = _RAND_5542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5543 = {1{`RANDOM}};
  _T_2982_re = _RAND_5543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5544 = {1{`RANDOM}};
  _T_2982_im = _RAND_5544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5545 = {1{`RANDOM}};
  _T_2983_re = _RAND_5545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5546 = {1{`RANDOM}};
  _T_2983_im = _RAND_5546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5547 = {1{`RANDOM}};
  _T_2984_re = _RAND_5547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5548 = {1{`RANDOM}};
  _T_2984_im = _RAND_5548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5549 = {1{`RANDOM}};
  _T_2985_re = _RAND_5549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5550 = {1{`RANDOM}};
  _T_2985_im = _RAND_5550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5551 = {1{`RANDOM}};
  _T_2986_re = _RAND_5551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5552 = {1{`RANDOM}};
  _T_2986_im = _RAND_5552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5553 = {1{`RANDOM}};
  _T_2987_re = _RAND_5553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5554 = {1{`RANDOM}};
  _T_2987_im = _RAND_5554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5555 = {1{`RANDOM}};
  _T_2988_re = _RAND_5555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5556 = {1{`RANDOM}};
  _T_2988_im = _RAND_5556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5557 = {1{`RANDOM}};
  _T_2989_re = _RAND_5557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5558 = {1{`RANDOM}};
  _T_2989_im = _RAND_5558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5559 = {1{`RANDOM}};
  _T_2990_re = _RAND_5559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5560 = {1{`RANDOM}};
  _T_2990_im = _RAND_5560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5561 = {1{`RANDOM}};
  _T_2991_re = _RAND_5561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5562 = {1{`RANDOM}};
  _T_2991_im = _RAND_5562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5563 = {1{`RANDOM}};
  _T_2992_re = _RAND_5563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5564 = {1{`RANDOM}};
  _T_2992_im = _RAND_5564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5565 = {1{`RANDOM}};
  _T_2993_re = _RAND_5565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5566 = {1{`RANDOM}};
  _T_2993_im = _RAND_5566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5567 = {1{`RANDOM}};
  _T_2994_re = _RAND_5567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5568 = {1{`RANDOM}};
  _T_2994_im = _RAND_5568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5569 = {1{`RANDOM}};
  _T_2995_re = _RAND_5569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5570 = {1{`RANDOM}};
  _T_2995_im = _RAND_5570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5571 = {1{`RANDOM}};
  _T_2996_re = _RAND_5571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5572 = {1{`RANDOM}};
  _T_2996_im = _RAND_5572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5573 = {1{`RANDOM}};
  _T_2997_re = _RAND_5573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5574 = {1{`RANDOM}};
  _T_2997_im = _RAND_5574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5575 = {1{`RANDOM}};
  _T_2998_re = _RAND_5575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5576 = {1{`RANDOM}};
  _T_2998_im = _RAND_5576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5577 = {1{`RANDOM}};
  _T_2999_re = _RAND_5577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5578 = {1{`RANDOM}};
  _T_2999_im = _RAND_5578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5579 = {1{`RANDOM}};
  _T_3000_re = _RAND_5579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5580 = {1{`RANDOM}};
  _T_3000_im = _RAND_5580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5581 = {1{`RANDOM}};
  _T_3001_re = _RAND_5581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5582 = {1{`RANDOM}};
  _T_3001_im = _RAND_5582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5583 = {1{`RANDOM}};
  _T_3002_re = _RAND_5583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5584 = {1{`RANDOM}};
  _T_3002_im = _RAND_5584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5585 = {1{`RANDOM}};
  _T_3003_re = _RAND_5585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5586 = {1{`RANDOM}};
  _T_3003_im = _RAND_5586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5587 = {1{`RANDOM}};
  _T_3004_re = _RAND_5587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5588 = {1{`RANDOM}};
  _T_3004_im = _RAND_5588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5589 = {1{`RANDOM}};
  _T_3005_re = _RAND_5589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5590 = {1{`RANDOM}};
  _T_3005_im = _RAND_5590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5591 = {1{`RANDOM}};
  _T_3006_re = _RAND_5591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5592 = {1{`RANDOM}};
  _T_3006_im = _RAND_5592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5593 = {1{`RANDOM}};
  _T_3007_re = _RAND_5593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5594 = {1{`RANDOM}};
  _T_3007_im = _RAND_5594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5595 = {1{`RANDOM}};
  _T_3008_re = _RAND_5595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5596 = {1{`RANDOM}};
  _T_3008_im = _RAND_5596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5597 = {1{`RANDOM}};
  _T_3009_re = _RAND_5597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5598 = {1{`RANDOM}};
  _T_3009_im = _RAND_5598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5599 = {1{`RANDOM}};
  _T_3010_re = _RAND_5599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5600 = {1{`RANDOM}};
  _T_3010_im = _RAND_5600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5601 = {1{`RANDOM}};
  _T_3011_re = _RAND_5601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5602 = {1{`RANDOM}};
  _T_3011_im = _RAND_5602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5603 = {1{`RANDOM}};
  _T_3012_re = _RAND_5603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5604 = {1{`RANDOM}};
  _T_3012_im = _RAND_5604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5605 = {1{`RANDOM}};
  _T_3013_re = _RAND_5605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5606 = {1{`RANDOM}};
  _T_3013_im = _RAND_5606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5607 = {1{`RANDOM}};
  _T_3014_re = _RAND_5607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5608 = {1{`RANDOM}};
  _T_3014_im = _RAND_5608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5609 = {1{`RANDOM}};
  _T_3015_re = _RAND_5609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5610 = {1{`RANDOM}};
  _T_3015_im = _RAND_5610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5611 = {1{`RANDOM}};
  _T_3016_re = _RAND_5611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5612 = {1{`RANDOM}};
  _T_3016_im = _RAND_5612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5613 = {1{`RANDOM}};
  _T_3017_re = _RAND_5613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5614 = {1{`RANDOM}};
  _T_3017_im = _RAND_5614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5615 = {1{`RANDOM}};
  _T_3018_re = _RAND_5615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5616 = {1{`RANDOM}};
  _T_3018_im = _RAND_5616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5617 = {1{`RANDOM}};
  _T_3019_re = _RAND_5617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5618 = {1{`RANDOM}};
  _T_3019_im = _RAND_5618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5619 = {1{`RANDOM}};
  _T_3020_re = _RAND_5619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5620 = {1{`RANDOM}};
  _T_3020_im = _RAND_5620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5621 = {1{`RANDOM}};
  _T_3021_re = _RAND_5621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5622 = {1{`RANDOM}};
  _T_3021_im = _RAND_5622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5623 = {1{`RANDOM}};
  _T_3022_re = _RAND_5623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5624 = {1{`RANDOM}};
  _T_3022_im = _RAND_5624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5625 = {1{`RANDOM}};
  _T_3023_re = _RAND_5625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5626 = {1{`RANDOM}};
  _T_3023_im = _RAND_5626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5627 = {1{`RANDOM}};
  _T_3024_re = _RAND_5627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5628 = {1{`RANDOM}};
  _T_3024_im = _RAND_5628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5629 = {1{`RANDOM}};
  _T_3025_re = _RAND_5629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5630 = {1{`RANDOM}};
  _T_3025_im = _RAND_5630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5631 = {1{`RANDOM}};
  _T_3026_re = _RAND_5631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5632 = {1{`RANDOM}};
  _T_3026_im = _RAND_5632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5633 = {1{`RANDOM}};
  _T_3027_re = _RAND_5633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5634 = {1{`RANDOM}};
  _T_3027_im = _RAND_5634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5635 = {1{`RANDOM}};
  _T_3028_re = _RAND_5635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5636 = {1{`RANDOM}};
  _T_3028_im = _RAND_5636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5637 = {1{`RANDOM}};
  _T_3029_re = _RAND_5637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5638 = {1{`RANDOM}};
  _T_3029_im = _RAND_5638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5639 = {1{`RANDOM}};
  _T_3032_re = _RAND_5639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5640 = {1{`RANDOM}};
  _T_3032_im = _RAND_5640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5641 = {1{`RANDOM}};
  _T_3033_re = _RAND_5641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5642 = {1{`RANDOM}};
  _T_3033_im = _RAND_5642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5643 = {1{`RANDOM}};
  _T_3034_re = _RAND_5643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5644 = {1{`RANDOM}};
  _T_3034_im = _RAND_5644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5645 = {1{`RANDOM}};
  _T_3035_re = _RAND_5645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5646 = {1{`RANDOM}};
  _T_3035_im = _RAND_5646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5647 = {1{`RANDOM}};
  _T_3036_re = _RAND_5647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5648 = {1{`RANDOM}};
  _T_3036_im = _RAND_5648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5649 = {1{`RANDOM}};
  _T_3037_re = _RAND_5649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5650 = {1{`RANDOM}};
  _T_3037_im = _RAND_5650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5651 = {1{`RANDOM}};
  _T_3038_re = _RAND_5651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5652 = {1{`RANDOM}};
  _T_3038_im = _RAND_5652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5653 = {1{`RANDOM}};
  _T_3039_re = _RAND_5653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5654 = {1{`RANDOM}};
  _T_3039_im = _RAND_5654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5655 = {1{`RANDOM}};
  _T_3040_re = _RAND_5655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5656 = {1{`RANDOM}};
  _T_3040_im = _RAND_5656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5657 = {1{`RANDOM}};
  _T_3041_re = _RAND_5657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5658 = {1{`RANDOM}};
  _T_3041_im = _RAND_5658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5659 = {1{`RANDOM}};
  _T_3042_re = _RAND_5659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5660 = {1{`RANDOM}};
  _T_3042_im = _RAND_5660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5661 = {1{`RANDOM}};
  _T_3043_re = _RAND_5661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5662 = {1{`RANDOM}};
  _T_3043_im = _RAND_5662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5663 = {1{`RANDOM}};
  _T_3044_re = _RAND_5663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5664 = {1{`RANDOM}};
  _T_3044_im = _RAND_5664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5665 = {1{`RANDOM}};
  _T_3045_re = _RAND_5665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5666 = {1{`RANDOM}};
  _T_3045_im = _RAND_5666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5667 = {1{`RANDOM}};
  _T_3046_re = _RAND_5667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5668 = {1{`RANDOM}};
  _T_3046_im = _RAND_5668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5669 = {1{`RANDOM}};
  _T_3047_re = _RAND_5669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5670 = {1{`RANDOM}};
  _T_3047_im = _RAND_5670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5671 = {1{`RANDOM}};
  _T_3048_re = _RAND_5671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5672 = {1{`RANDOM}};
  _T_3048_im = _RAND_5672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5673 = {1{`RANDOM}};
  _T_3049_re = _RAND_5673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5674 = {1{`RANDOM}};
  _T_3049_im = _RAND_5674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5675 = {1{`RANDOM}};
  _T_3050_re = _RAND_5675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5676 = {1{`RANDOM}};
  _T_3050_im = _RAND_5676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5677 = {1{`RANDOM}};
  _T_3051_re = _RAND_5677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5678 = {1{`RANDOM}};
  _T_3051_im = _RAND_5678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5679 = {1{`RANDOM}};
  _T_3052_re = _RAND_5679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5680 = {1{`RANDOM}};
  _T_3052_im = _RAND_5680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5681 = {1{`RANDOM}};
  _T_3053_re = _RAND_5681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5682 = {1{`RANDOM}};
  _T_3053_im = _RAND_5682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5683 = {1{`RANDOM}};
  _T_3054_re = _RAND_5683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5684 = {1{`RANDOM}};
  _T_3054_im = _RAND_5684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5685 = {1{`RANDOM}};
  _T_3055_re = _RAND_5685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5686 = {1{`RANDOM}};
  _T_3055_im = _RAND_5686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5687 = {1{`RANDOM}};
  _T_3056_re = _RAND_5687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5688 = {1{`RANDOM}};
  _T_3056_im = _RAND_5688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5689 = {1{`RANDOM}};
  _T_3057_re = _RAND_5689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5690 = {1{`RANDOM}};
  _T_3057_im = _RAND_5690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5691 = {1{`RANDOM}};
  _T_3058_re = _RAND_5691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5692 = {1{`RANDOM}};
  _T_3058_im = _RAND_5692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5693 = {1{`RANDOM}};
  _T_3059_re = _RAND_5693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5694 = {1{`RANDOM}};
  _T_3059_im = _RAND_5694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5695 = {1{`RANDOM}};
  _T_3060_re = _RAND_5695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5696 = {1{`RANDOM}};
  _T_3060_im = _RAND_5696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5697 = {1{`RANDOM}};
  _T_3061_re = _RAND_5697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5698 = {1{`RANDOM}};
  _T_3061_im = _RAND_5698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5699 = {1{`RANDOM}};
  _T_3062_re = _RAND_5699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5700 = {1{`RANDOM}};
  _T_3062_im = _RAND_5700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5701 = {1{`RANDOM}};
  _T_3063_re = _RAND_5701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5702 = {1{`RANDOM}};
  _T_3063_im = _RAND_5702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5703 = {1{`RANDOM}};
  _T_3064_re = _RAND_5703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5704 = {1{`RANDOM}};
  _T_3064_im = _RAND_5704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5705 = {1{`RANDOM}};
  _T_3065_re = _RAND_5705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5706 = {1{`RANDOM}};
  _T_3065_im = _RAND_5706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5707 = {1{`RANDOM}};
  _T_3066_re = _RAND_5707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5708 = {1{`RANDOM}};
  _T_3066_im = _RAND_5708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5709 = {1{`RANDOM}};
  _T_3067_re = _RAND_5709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5710 = {1{`RANDOM}};
  _T_3067_im = _RAND_5710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5711 = {1{`RANDOM}};
  _T_3068_re = _RAND_5711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5712 = {1{`RANDOM}};
  _T_3068_im = _RAND_5712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5713 = {1{`RANDOM}};
  _T_3069_re = _RAND_5713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5714 = {1{`RANDOM}};
  _T_3069_im = _RAND_5714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5715 = {1{`RANDOM}};
  _T_3070_re = _RAND_5715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5716 = {1{`RANDOM}};
  _T_3070_im = _RAND_5716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5717 = {1{`RANDOM}};
  _T_3071_re = _RAND_5717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5718 = {1{`RANDOM}};
  _T_3071_im = _RAND_5718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5719 = {1{`RANDOM}};
  _T_3072_re = _RAND_5719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5720 = {1{`RANDOM}};
  _T_3072_im = _RAND_5720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5721 = {1{`RANDOM}};
  _T_3073_re = _RAND_5721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5722 = {1{`RANDOM}};
  _T_3073_im = _RAND_5722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5723 = {1{`RANDOM}};
  _T_3074_re = _RAND_5723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5724 = {1{`RANDOM}};
  _T_3074_im = _RAND_5724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5725 = {1{`RANDOM}};
  _T_3075_re = _RAND_5725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5726 = {1{`RANDOM}};
  _T_3075_im = _RAND_5726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5727 = {1{`RANDOM}};
  _T_3076_re = _RAND_5727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5728 = {1{`RANDOM}};
  _T_3076_im = _RAND_5728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5729 = {1{`RANDOM}};
  _T_3077_re = _RAND_5729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5730 = {1{`RANDOM}};
  _T_3077_im = _RAND_5730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5731 = {1{`RANDOM}};
  _T_3078_re = _RAND_5731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5732 = {1{`RANDOM}};
  _T_3078_im = _RAND_5732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5733 = {1{`RANDOM}};
  _T_3079_re = _RAND_5733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5734 = {1{`RANDOM}};
  _T_3079_im = _RAND_5734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5735 = {1{`RANDOM}};
  _T_3080_re = _RAND_5735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5736 = {1{`RANDOM}};
  _T_3080_im = _RAND_5736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5737 = {1{`RANDOM}};
  _T_3081_re = _RAND_5737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5738 = {1{`RANDOM}};
  _T_3081_im = _RAND_5738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5739 = {1{`RANDOM}};
  _T_3082_re = _RAND_5739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5740 = {1{`RANDOM}};
  _T_3082_im = _RAND_5740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5741 = {1{`RANDOM}};
  _T_3083_re = _RAND_5741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5742 = {1{`RANDOM}};
  _T_3083_im = _RAND_5742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5743 = {1{`RANDOM}};
  _T_3084_re = _RAND_5743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5744 = {1{`RANDOM}};
  _T_3084_im = _RAND_5744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5745 = {1{`RANDOM}};
  _T_3085_re = _RAND_5745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5746 = {1{`RANDOM}};
  _T_3085_im = _RAND_5746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5747 = {1{`RANDOM}};
  _T_3086_re = _RAND_5747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5748 = {1{`RANDOM}};
  _T_3086_im = _RAND_5748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5749 = {1{`RANDOM}};
  _T_3087_re = _RAND_5749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5750 = {1{`RANDOM}};
  _T_3087_im = _RAND_5750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5751 = {1{`RANDOM}};
  _T_3088_re = _RAND_5751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5752 = {1{`RANDOM}};
  _T_3088_im = _RAND_5752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5753 = {1{`RANDOM}};
  _T_3089_re = _RAND_5753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5754 = {1{`RANDOM}};
  _T_3089_im = _RAND_5754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5755 = {1{`RANDOM}};
  _T_3090_re = _RAND_5755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5756 = {1{`RANDOM}};
  _T_3090_im = _RAND_5756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5757 = {1{`RANDOM}};
  _T_3091_re = _RAND_5757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5758 = {1{`RANDOM}};
  _T_3091_im = _RAND_5758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5759 = {1{`RANDOM}};
  _T_3092_re = _RAND_5759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5760 = {1{`RANDOM}};
  _T_3092_im = _RAND_5760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5761 = {1{`RANDOM}};
  _T_3093_re = _RAND_5761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5762 = {1{`RANDOM}};
  _T_3093_im = _RAND_5762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5763 = {1{`RANDOM}};
  _T_3094_re = _RAND_5763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5764 = {1{`RANDOM}};
  _T_3094_im = _RAND_5764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5765 = {1{`RANDOM}};
  _T_3095_re = _RAND_5765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5766 = {1{`RANDOM}};
  _T_3095_im = _RAND_5766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5767 = {1{`RANDOM}};
  _T_3105_re = _RAND_5767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5768 = {1{`RANDOM}};
  _T_3105_im = _RAND_5768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5769 = {1{`RANDOM}};
  _T_3106_re = _RAND_5769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5770 = {1{`RANDOM}};
  _T_3106_im = _RAND_5770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5771 = {1{`RANDOM}};
  _T_3107_re = _RAND_5771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5772 = {1{`RANDOM}};
  _T_3107_im = _RAND_5772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5773 = {1{`RANDOM}};
  _T_3108_re = _RAND_5773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5774 = {1{`RANDOM}};
  _T_3108_im = _RAND_5774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5775 = {1{`RANDOM}};
  _T_3109_re = _RAND_5775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5776 = {1{`RANDOM}};
  _T_3109_im = _RAND_5776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5777 = {1{`RANDOM}};
  _T_3110_re = _RAND_5777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5778 = {1{`RANDOM}};
  _T_3110_im = _RAND_5778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5779 = {1{`RANDOM}};
  _T_3111_re = _RAND_5779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5780 = {1{`RANDOM}};
  _T_3111_im = _RAND_5780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5781 = {1{`RANDOM}};
  _T_3112_re = _RAND_5781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5782 = {1{`RANDOM}};
  _T_3112_im = _RAND_5782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5783 = {1{`RANDOM}};
  _T_3113_re = _RAND_5783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5784 = {1{`RANDOM}};
  _T_3113_im = _RAND_5784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5785 = {1{`RANDOM}};
  _T_3114_re = _RAND_5785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5786 = {1{`RANDOM}};
  _T_3114_im = _RAND_5786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5787 = {1{`RANDOM}};
  _T_3115_re = _RAND_5787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5788 = {1{`RANDOM}};
  _T_3115_im = _RAND_5788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5789 = {1{`RANDOM}};
  _T_3116_re = _RAND_5789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5790 = {1{`RANDOM}};
  _T_3116_im = _RAND_5790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5791 = {1{`RANDOM}};
  _T_3117_re = _RAND_5791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5792 = {1{`RANDOM}};
  _T_3117_im = _RAND_5792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5793 = {1{`RANDOM}};
  _T_3118_re = _RAND_5793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5794 = {1{`RANDOM}};
  _T_3118_im = _RAND_5794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5795 = {1{`RANDOM}};
  _T_3119_re = _RAND_5795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5796 = {1{`RANDOM}};
  _T_3119_im = _RAND_5796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5797 = {1{`RANDOM}};
  _T_3120_re = _RAND_5797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5798 = {1{`RANDOM}};
  _T_3120_im = _RAND_5798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5799 = {1{`RANDOM}};
  _T_3121_re = _RAND_5799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5800 = {1{`RANDOM}};
  _T_3121_im = _RAND_5800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5801 = {1{`RANDOM}};
  _T_3122_re = _RAND_5801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5802 = {1{`RANDOM}};
  _T_3122_im = _RAND_5802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5803 = {1{`RANDOM}};
  _T_3123_re = _RAND_5803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5804 = {1{`RANDOM}};
  _T_3123_im = _RAND_5804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5805 = {1{`RANDOM}};
  _T_3124_re = _RAND_5805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5806 = {1{`RANDOM}};
  _T_3124_im = _RAND_5806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5807 = {1{`RANDOM}};
  _T_3125_re = _RAND_5807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5808 = {1{`RANDOM}};
  _T_3125_im = _RAND_5808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5809 = {1{`RANDOM}};
  _T_3126_re = _RAND_5809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5810 = {1{`RANDOM}};
  _T_3126_im = _RAND_5810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5811 = {1{`RANDOM}};
  _T_3127_re = _RAND_5811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5812 = {1{`RANDOM}};
  _T_3127_im = _RAND_5812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5813 = {1{`RANDOM}};
  _T_3128_re = _RAND_5813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5814 = {1{`RANDOM}};
  _T_3128_im = _RAND_5814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5815 = {1{`RANDOM}};
  _T_3129_re = _RAND_5815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5816 = {1{`RANDOM}};
  _T_3129_im = _RAND_5816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5817 = {1{`RANDOM}};
  _T_3130_re = _RAND_5817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5818 = {1{`RANDOM}};
  _T_3130_im = _RAND_5818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5819 = {1{`RANDOM}};
  _T_3131_re = _RAND_5819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5820 = {1{`RANDOM}};
  _T_3131_im = _RAND_5820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5821 = {1{`RANDOM}};
  _T_3132_re = _RAND_5821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5822 = {1{`RANDOM}};
  _T_3132_im = _RAND_5822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5823 = {1{`RANDOM}};
  _T_3133_re = _RAND_5823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5824 = {1{`RANDOM}};
  _T_3133_im = _RAND_5824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5825 = {1{`RANDOM}};
  _T_3134_re = _RAND_5825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5826 = {1{`RANDOM}};
  _T_3134_im = _RAND_5826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5827 = {1{`RANDOM}};
  _T_3135_re = _RAND_5827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5828 = {1{`RANDOM}};
  _T_3135_im = _RAND_5828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5829 = {1{`RANDOM}};
  _T_3136_re = _RAND_5829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5830 = {1{`RANDOM}};
  _T_3136_im = _RAND_5830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5831 = {1{`RANDOM}};
  _T_3137_re = _RAND_5831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5832 = {1{`RANDOM}};
  _T_3137_im = _RAND_5832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5833 = {1{`RANDOM}};
  _T_3138_re = _RAND_5833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5834 = {1{`RANDOM}};
  _T_3138_im = _RAND_5834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5835 = {1{`RANDOM}};
  _T_3139_re = _RAND_5835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5836 = {1{`RANDOM}};
  _T_3139_im = _RAND_5836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5837 = {1{`RANDOM}};
  _T_3140_re = _RAND_5837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5838 = {1{`RANDOM}};
  _T_3140_im = _RAND_5838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5839 = {1{`RANDOM}};
  _T_3141_re = _RAND_5839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5840 = {1{`RANDOM}};
  _T_3141_im = _RAND_5840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5841 = {1{`RANDOM}};
  _T_3142_re = _RAND_5841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5842 = {1{`RANDOM}};
  _T_3142_im = _RAND_5842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5843 = {1{`RANDOM}};
  _T_3143_re = _RAND_5843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5844 = {1{`RANDOM}};
  _T_3143_im = _RAND_5844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5845 = {1{`RANDOM}};
  _T_3144_re = _RAND_5845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5846 = {1{`RANDOM}};
  _T_3144_im = _RAND_5846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5847 = {1{`RANDOM}};
  _T_3145_re = _RAND_5847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5848 = {1{`RANDOM}};
  _T_3145_im = _RAND_5848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5849 = {1{`RANDOM}};
  _T_3146_re = _RAND_5849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5850 = {1{`RANDOM}};
  _T_3146_im = _RAND_5850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5851 = {1{`RANDOM}};
  _T_3147_re = _RAND_5851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5852 = {1{`RANDOM}};
  _T_3147_im = _RAND_5852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5853 = {1{`RANDOM}};
  _T_3148_re = _RAND_5853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5854 = {1{`RANDOM}};
  _T_3148_im = _RAND_5854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5855 = {1{`RANDOM}};
  _T_3149_re = _RAND_5855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5856 = {1{`RANDOM}};
  _T_3149_im = _RAND_5856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5857 = {1{`RANDOM}};
  _T_3150_re = _RAND_5857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5858 = {1{`RANDOM}};
  _T_3150_im = _RAND_5858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5859 = {1{`RANDOM}};
  _T_3151_re = _RAND_5859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5860 = {1{`RANDOM}};
  _T_3151_im = _RAND_5860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5861 = {1{`RANDOM}};
  _T_3152_re = _RAND_5861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5862 = {1{`RANDOM}};
  _T_3152_im = _RAND_5862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5863 = {1{`RANDOM}};
  _T_3153_re = _RAND_5863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5864 = {1{`RANDOM}};
  _T_3153_im = _RAND_5864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5865 = {1{`RANDOM}};
  _T_3154_re = _RAND_5865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5866 = {1{`RANDOM}};
  _T_3154_im = _RAND_5866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5867 = {1{`RANDOM}};
  _T_3155_re = _RAND_5867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5868 = {1{`RANDOM}};
  _T_3155_im = _RAND_5868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5869 = {1{`RANDOM}};
  _T_3156_re = _RAND_5869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5870 = {1{`RANDOM}};
  _T_3156_im = _RAND_5870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5871 = {1{`RANDOM}};
  _T_3157_re = _RAND_5871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5872 = {1{`RANDOM}};
  _T_3157_im = _RAND_5872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5873 = {1{`RANDOM}};
  _T_3158_re = _RAND_5873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5874 = {1{`RANDOM}};
  _T_3158_im = _RAND_5874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5875 = {1{`RANDOM}};
  _T_3159_re = _RAND_5875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5876 = {1{`RANDOM}};
  _T_3159_im = _RAND_5876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5877 = {1{`RANDOM}};
  _T_3160_re = _RAND_5877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5878 = {1{`RANDOM}};
  _T_3160_im = _RAND_5878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5879 = {1{`RANDOM}};
  _T_3161_re = _RAND_5879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5880 = {1{`RANDOM}};
  _T_3161_im = _RAND_5880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5881 = {1{`RANDOM}};
  _T_3162_re = _RAND_5881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5882 = {1{`RANDOM}};
  _T_3162_im = _RAND_5882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5883 = {1{`RANDOM}};
  _T_3163_re = _RAND_5883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5884 = {1{`RANDOM}};
  _T_3163_im = _RAND_5884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5885 = {1{`RANDOM}};
  _T_3164_re = _RAND_5885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5886 = {1{`RANDOM}};
  _T_3164_im = _RAND_5886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5887 = {1{`RANDOM}};
  _T_3165_re = _RAND_5887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5888 = {1{`RANDOM}};
  _T_3165_im = _RAND_5888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5889 = {1{`RANDOM}};
  _T_3166_re = _RAND_5889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5890 = {1{`RANDOM}};
  _T_3166_im = _RAND_5890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5891 = {1{`RANDOM}};
  _T_3167_re = _RAND_5891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5892 = {1{`RANDOM}};
  _T_3167_im = _RAND_5892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5893 = {1{`RANDOM}};
  _T_3168_re = _RAND_5893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5894 = {1{`RANDOM}};
  _T_3168_im = _RAND_5894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5895 = {1{`RANDOM}};
  _T_3171_re = _RAND_5895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5896 = {1{`RANDOM}};
  _T_3171_im = _RAND_5896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5897 = {1{`RANDOM}};
  _T_3172_re = _RAND_5897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5898 = {1{`RANDOM}};
  _T_3172_im = _RAND_5898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5899 = {1{`RANDOM}};
  _T_3173_re = _RAND_5899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5900 = {1{`RANDOM}};
  _T_3173_im = _RAND_5900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5901 = {1{`RANDOM}};
  _T_3174_re = _RAND_5901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5902 = {1{`RANDOM}};
  _T_3174_im = _RAND_5902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5903 = {1{`RANDOM}};
  _T_3175_re = _RAND_5903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5904 = {1{`RANDOM}};
  _T_3175_im = _RAND_5904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5905 = {1{`RANDOM}};
  _T_3176_re = _RAND_5905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5906 = {1{`RANDOM}};
  _T_3176_im = _RAND_5906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5907 = {1{`RANDOM}};
  _T_3177_re = _RAND_5907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5908 = {1{`RANDOM}};
  _T_3177_im = _RAND_5908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5909 = {1{`RANDOM}};
  _T_3178_re = _RAND_5909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5910 = {1{`RANDOM}};
  _T_3178_im = _RAND_5910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5911 = {1{`RANDOM}};
  _T_3179_re = _RAND_5911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5912 = {1{`RANDOM}};
  _T_3179_im = _RAND_5912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5913 = {1{`RANDOM}};
  _T_3180_re = _RAND_5913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5914 = {1{`RANDOM}};
  _T_3180_im = _RAND_5914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5915 = {1{`RANDOM}};
  _T_3181_re = _RAND_5915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5916 = {1{`RANDOM}};
  _T_3181_im = _RAND_5916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5917 = {1{`RANDOM}};
  _T_3182_re = _RAND_5917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5918 = {1{`RANDOM}};
  _T_3182_im = _RAND_5918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5919 = {1{`RANDOM}};
  _T_3183_re = _RAND_5919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5920 = {1{`RANDOM}};
  _T_3183_im = _RAND_5920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5921 = {1{`RANDOM}};
  _T_3184_re = _RAND_5921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5922 = {1{`RANDOM}};
  _T_3184_im = _RAND_5922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5923 = {1{`RANDOM}};
  _T_3185_re = _RAND_5923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5924 = {1{`RANDOM}};
  _T_3185_im = _RAND_5924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5925 = {1{`RANDOM}};
  _T_3186_re = _RAND_5925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5926 = {1{`RANDOM}};
  _T_3186_im = _RAND_5926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5927 = {1{`RANDOM}};
  _T_3187_re = _RAND_5927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5928 = {1{`RANDOM}};
  _T_3187_im = _RAND_5928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5929 = {1{`RANDOM}};
  _T_3188_re = _RAND_5929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5930 = {1{`RANDOM}};
  _T_3188_im = _RAND_5930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5931 = {1{`RANDOM}};
  _T_3189_re = _RAND_5931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5932 = {1{`RANDOM}};
  _T_3189_im = _RAND_5932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5933 = {1{`RANDOM}};
  _T_3190_re = _RAND_5933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5934 = {1{`RANDOM}};
  _T_3190_im = _RAND_5934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5935 = {1{`RANDOM}};
  _T_3191_re = _RAND_5935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5936 = {1{`RANDOM}};
  _T_3191_im = _RAND_5936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5937 = {1{`RANDOM}};
  _T_3192_re = _RAND_5937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5938 = {1{`RANDOM}};
  _T_3192_im = _RAND_5938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5939 = {1{`RANDOM}};
  _T_3193_re = _RAND_5939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5940 = {1{`RANDOM}};
  _T_3193_im = _RAND_5940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5941 = {1{`RANDOM}};
  _T_3194_re = _RAND_5941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5942 = {1{`RANDOM}};
  _T_3194_im = _RAND_5942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5943 = {1{`RANDOM}};
  _T_3195_re = _RAND_5943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5944 = {1{`RANDOM}};
  _T_3195_im = _RAND_5944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5945 = {1{`RANDOM}};
  _T_3196_re = _RAND_5945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5946 = {1{`RANDOM}};
  _T_3196_im = _RAND_5946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5947 = {1{`RANDOM}};
  _T_3197_re = _RAND_5947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5948 = {1{`RANDOM}};
  _T_3197_im = _RAND_5948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5949 = {1{`RANDOM}};
  _T_3198_re = _RAND_5949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5950 = {1{`RANDOM}};
  _T_3198_im = _RAND_5950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5951 = {1{`RANDOM}};
  _T_3199_re = _RAND_5951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5952 = {1{`RANDOM}};
  _T_3199_im = _RAND_5952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5953 = {1{`RANDOM}};
  _T_3200_re = _RAND_5953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5954 = {1{`RANDOM}};
  _T_3200_im = _RAND_5954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5955 = {1{`RANDOM}};
  _T_3201_re = _RAND_5955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5956 = {1{`RANDOM}};
  _T_3201_im = _RAND_5956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5957 = {1{`RANDOM}};
  _T_3202_re = _RAND_5957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5958 = {1{`RANDOM}};
  _T_3202_im = _RAND_5958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5959 = {1{`RANDOM}};
  _T_3212_re = _RAND_5959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5960 = {1{`RANDOM}};
  _T_3212_im = _RAND_5960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5961 = {1{`RANDOM}};
  _T_3213_re = _RAND_5961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5962 = {1{`RANDOM}};
  _T_3213_im = _RAND_5962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5963 = {1{`RANDOM}};
  _T_3214_re = _RAND_5963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5964 = {1{`RANDOM}};
  _T_3214_im = _RAND_5964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5965 = {1{`RANDOM}};
  _T_3215_re = _RAND_5965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5966 = {1{`RANDOM}};
  _T_3215_im = _RAND_5966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5967 = {1{`RANDOM}};
  _T_3216_re = _RAND_5967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5968 = {1{`RANDOM}};
  _T_3216_im = _RAND_5968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5969 = {1{`RANDOM}};
  _T_3217_re = _RAND_5969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5970 = {1{`RANDOM}};
  _T_3217_im = _RAND_5970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5971 = {1{`RANDOM}};
  _T_3218_re = _RAND_5971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5972 = {1{`RANDOM}};
  _T_3218_im = _RAND_5972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5973 = {1{`RANDOM}};
  _T_3219_re = _RAND_5973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5974 = {1{`RANDOM}};
  _T_3219_im = _RAND_5974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5975 = {1{`RANDOM}};
  _T_3220_re = _RAND_5975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5976 = {1{`RANDOM}};
  _T_3220_im = _RAND_5976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5977 = {1{`RANDOM}};
  _T_3221_re = _RAND_5977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5978 = {1{`RANDOM}};
  _T_3221_im = _RAND_5978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5979 = {1{`RANDOM}};
  _T_3222_re = _RAND_5979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5980 = {1{`RANDOM}};
  _T_3222_im = _RAND_5980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5981 = {1{`RANDOM}};
  _T_3223_re = _RAND_5981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5982 = {1{`RANDOM}};
  _T_3223_im = _RAND_5982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5983 = {1{`RANDOM}};
  _T_3224_re = _RAND_5983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5984 = {1{`RANDOM}};
  _T_3224_im = _RAND_5984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5985 = {1{`RANDOM}};
  _T_3225_re = _RAND_5985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5986 = {1{`RANDOM}};
  _T_3225_im = _RAND_5986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5987 = {1{`RANDOM}};
  _T_3226_re = _RAND_5987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5988 = {1{`RANDOM}};
  _T_3226_im = _RAND_5988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5989 = {1{`RANDOM}};
  _T_3227_re = _RAND_5989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5990 = {1{`RANDOM}};
  _T_3227_im = _RAND_5990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5991 = {1{`RANDOM}};
  _T_3228_re = _RAND_5991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5992 = {1{`RANDOM}};
  _T_3228_im = _RAND_5992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5993 = {1{`RANDOM}};
  _T_3229_re = _RAND_5993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5994 = {1{`RANDOM}};
  _T_3229_im = _RAND_5994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5995 = {1{`RANDOM}};
  _T_3230_re = _RAND_5995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5996 = {1{`RANDOM}};
  _T_3230_im = _RAND_5996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5997 = {1{`RANDOM}};
  _T_3231_re = _RAND_5997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5998 = {1{`RANDOM}};
  _T_3231_im = _RAND_5998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5999 = {1{`RANDOM}};
  _T_3232_re = _RAND_5999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6000 = {1{`RANDOM}};
  _T_3232_im = _RAND_6000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6001 = {1{`RANDOM}};
  _T_3233_re = _RAND_6001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6002 = {1{`RANDOM}};
  _T_3233_im = _RAND_6002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6003 = {1{`RANDOM}};
  _T_3234_re = _RAND_6003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6004 = {1{`RANDOM}};
  _T_3234_im = _RAND_6004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6005 = {1{`RANDOM}};
  _T_3235_re = _RAND_6005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6006 = {1{`RANDOM}};
  _T_3235_im = _RAND_6006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6007 = {1{`RANDOM}};
  _T_3236_re = _RAND_6007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6008 = {1{`RANDOM}};
  _T_3236_im = _RAND_6008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6009 = {1{`RANDOM}};
  _T_3237_re = _RAND_6009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6010 = {1{`RANDOM}};
  _T_3237_im = _RAND_6010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6011 = {1{`RANDOM}};
  _T_3238_re = _RAND_6011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6012 = {1{`RANDOM}};
  _T_3238_im = _RAND_6012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6013 = {1{`RANDOM}};
  _T_3239_re = _RAND_6013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6014 = {1{`RANDOM}};
  _T_3239_im = _RAND_6014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6015 = {1{`RANDOM}};
  _T_3240_re = _RAND_6015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6016 = {1{`RANDOM}};
  _T_3240_im = _RAND_6016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6017 = {1{`RANDOM}};
  _T_3241_re = _RAND_6017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6018 = {1{`RANDOM}};
  _T_3241_im = _RAND_6018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6019 = {1{`RANDOM}};
  _T_3242_re = _RAND_6019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6020 = {1{`RANDOM}};
  _T_3242_im = _RAND_6020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6021 = {1{`RANDOM}};
  _T_3243_re = _RAND_6021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6022 = {1{`RANDOM}};
  _T_3243_im = _RAND_6022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6023 = {1{`RANDOM}};
  _T_3246_re = _RAND_6023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6024 = {1{`RANDOM}};
  _T_3246_im = _RAND_6024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6025 = {1{`RANDOM}};
  _T_3247_re = _RAND_6025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6026 = {1{`RANDOM}};
  _T_3247_im = _RAND_6026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6027 = {1{`RANDOM}};
  _T_3248_re = _RAND_6027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6028 = {1{`RANDOM}};
  _T_3248_im = _RAND_6028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6029 = {1{`RANDOM}};
  _T_3249_re = _RAND_6029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6030 = {1{`RANDOM}};
  _T_3249_im = _RAND_6030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6031 = {1{`RANDOM}};
  _T_3250_re = _RAND_6031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6032 = {1{`RANDOM}};
  _T_3250_im = _RAND_6032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6033 = {1{`RANDOM}};
  _T_3251_re = _RAND_6033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6034 = {1{`RANDOM}};
  _T_3251_im = _RAND_6034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6035 = {1{`RANDOM}};
  _T_3252_re = _RAND_6035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6036 = {1{`RANDOM}};
  _T_3252_im = _RAND_6036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6037 = {1{`RANDOM}};
  _T_3253_re = _RAND_6037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6038 = {1{`RANDOM}};
  _T_3253_im = _RAND_6038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6039 = {1{`RANDOM}};
  _T_3254_re = _RAND_6039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6040 = {1{`RANDOM}};
  _T_3254_im = _RAND_6040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6041 = {1{`RANDOM}};
  _T_3255_re = _RAND_6041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6042 = {1{`RANDOM}};
  _T_3255_im = _RAND_6042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6043 = {1{`RANDOM}};
  _T_3256_re = _RAND_6043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6044 = {1{`RANDOM}};
  _T_3256_im = _RAND_6044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6045 = {1{`RANDOM}};
  _T_3257_re = _RAND_6045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6046 = {1{`RANDOM}};
  _T_3257_im = _RAND_6046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6047 = {1{`RANDOM}};
  _T_3258_re = _RAND_6047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6048 = {1{`RANDOM}};
  _T_3258_im = _RAND_6048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6049 = {1{`RANDOM}};
  _T_3259_re = _RAND_6049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6050 = {1{`RANDOM}};
  _T_3259_im = _RAND_6050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6051 = {1{`RANDOM}};
  _T_3260_re = _RAND_6051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6052 = {1{`RANDOM}};
  _T_3260_im = _RAND_6052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6053 = {1{`RANDOM}};
  _T_3261_re = _RAND_6053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6054 = {1{`RANDOM}};
  _T_3261_im = _RAND_6054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6055 = {1{`RANDOM}};
  _T_3267_re = _RAND_6055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6056 = {1{`RANDOM}};
  _T_3267_im = _RAND_6056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6057 = {1{`RANDOM}};
  _T_3268_re = _RAND_6057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6058 = {1{`RANDOM}};
  _T_3268_im = _RAND_6058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6059 = {1{`RANDOM}};
  _T_3269_re = _RAND_6059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6060 = {1{`RANDOM}};
  _T_3269_im = _RAND_6060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6061 = {1{`RANDOM}};
  _T_3270_re = _RAND_6061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6062 = {1{`RANDOM}};
  _T_3270_im = _RAND_6062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6063 = {1{`RANDOM}};
  _T_3271_re = _RAND_6063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6064 = {1{`RANDOM}};
  _T_3271_im = _RAND_6064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6065 = {1{`RANDOM}};
  _T_3272_re = _RAND_6065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6066 = {1{`RANDOM}};
  _T_3272_im = _RAND_6066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6067 = {1{`RANDOM}};
  _T_3273_re = _RAND_6067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6068 = {1{`RANDOM}};
  _T_3273_im = _RAND_6068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6069 = {1{`RANDOM}};
  _T_3274_re = _RAND_6069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6070 = {1{`RANDOM}};
  _T_3274_im = _RAND_6070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6071 = {1{`RANDOM}};
  _T_3275_re = _RAND_6071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6072 = {1{`RANDOM}};
  _T_3275_im = _RAND_6072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6073 = {1{`RANDOM}};
  _T_3276_re = _RAND_6073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6074 = {1{`RANDOM}};
  _T_3276_im = _RAND_6074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6075 = {1{`RANDOM}};
  _T_3277_re = _RAND_6075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6076 = {1{`RANDOM}};
  _T_3277_im = _RAND_6076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6077 = {1{`RANDOM}};
  _T_3278_re = _RAND_6077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6078 = {1{`RANDOM}};
  _T_3278_im = _RAND_6078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6079 = {1{`RANDOM}};
  _T_3279_re = _RAND_6079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6080 = {1{`RANDOM}};
  _T_3279_im = _RAND_6080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6081 = {1{`RANDOM}};
  _T_3280_re = _RAND_6081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6082 = {1{`RANDOM}};
  _T_3280_im = _RAND_6082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6083 = {1{`RANDOM}};
  _T_3281_re = _RAND_6083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6084 = {1{`RANDOM}};
  _T_3281_im = _RAND_6084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6085 = {1{`RANDOM}};
  _T_3282_re = _RAND_6085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6086 = {1{`RANDOM}};
  _T_3282_im = _RAND_6086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6087 = {1{`RANDOM}};
  _T_3285_re = _RAND_6087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6088 = {1{`RANDOM}};
  _T_3285_im = _RAND_6088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6089 = {1{`RANDOM}};
  _T_3286_re = _RAND_6089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6090 = {1{`RANDOM}};
  _T_3286_im = _RAND_6090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6091 = {1{`RANDOM}};
  _T_3287_re = _RAND_6091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6092 = {1{`RANDOM}};
  _T_3287_im = _RAND_6092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6093 = {1{`RANDOM}};
  _T_3288_re = _RAND_6093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6094 = {1{`RANDOM}};
  _T_3288_im = _RAND_6094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6095 = {1{`RANDOM}};
  _T_3289_re = _RAND_6095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6096 = {1{`RANDOM}};
  _T_3289_im = _RAND_6096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6097 = {1{`RANDOM}};
  _T_3290_re = _RAND_6097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6098 = {1{`RANDOM}};
  _T_3290_im = _RAND_6098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6099 = {1{`RANDOM}};
  _T_3291_re = _RAND_6099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6100 = {1{`RANDOM}};
  _T_3291_im = _RAND_6100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6101 = {1{`RANDOM}};
  _T_3292_re = _RAND_6101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6102 = {1{`RANDOM}};
  _T_3292_im = _RAND_6102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6103 = {1{`RANDOM}};
  _T_3298_re = _RAND_6103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6104 = {1{`RANDOM}};
  _T_3298_im = _RAND_6104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6105 = {1{`RANDOM}};
  _T_3299_re = _RAND_6105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6106 = {1{`RANDOM}};
  _T_3299_im = _RAND_6106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6107 = {1{`RANDOM}};
  _T_3300_re = _RAND_6107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6108 = {1{`RANDOM}};
  _T_3300_im = _RAND_6108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6109 = {1{`RANDOM}};
  _T_3301_re = _RAND_6109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6110 = {1{`RANDOM}};
  _T_3301_im = _RAND_6110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6111 = {1{`RANDOM}};
  _T_3302_re = _RAND_6111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6112 = {1{`RANDOM}};
  _T_3302_im = _RAND_6112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6113 = {1{`RANDOM}};
  _T_3303_re = _RAND_6113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6114 = {1{`RANDOM}};
  _T_3303_im = _RAND_6114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6115 = {1{`RANDOM}};
  _T_3304_re = _RAND_6115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6116 = {1{`RANDOM}};
  _T_3304_im = _RAND_6116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6117 = {1{`RANDOM}};
  _T_3305_re = _RAND_6117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6118 = {1{`RANDOM}};
  _T_3305_im = _RAND_6118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6119 = {1{`RANDOM}};
  _T_3308_re = _RAND_6119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6120 = {1{`RANDOM}};
  _T_3308_im = _RAND_6120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6121 = {1{`RANDOM}};
  _T_3309_re = _RAND_6121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6122 = {1{`RANDOM}};
  _T_3309_im = _RAND_6122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6123 = {1{`RANDOM}};
  _T_3310_re = _RAND_6123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6124 = {1{`RANDOM}};
  _T_3310_im = _RAND_6124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6125 = {1{`RANDOM}};
  _T_3311_re = _RAND_6125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6126 = {1{`RANDOM}};
  _T_3311_im = _RAND_6126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6127 = {1{`RANDOM}};
  _T_3317_re = _RAND_6127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6128 = {1{`RANDOM}};
  _T_3317_im = _RAND_6128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6129 = {1{`RANDOM}};
  _T_3318_re = _RAND_6129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6130 = {1{`RANDOM}};
  _T_3318_im = _RAND_6130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6131 = {1{`RANDOM}};
  _T_3319_re = _RAND_6131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6132 = {1{`RANDOM}};
  _T_3319_im = _RAND_6132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6133 = {1{`RANDOM}};
  _T_3320_re = _RAND_6133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6134 = {1{`RANDOM}};
  _T_3320_im = _RAND_6134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6135 = {1{`RANDOM}};
  _T_3323_re = _RAND_6135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6136 = {1{`RANDOM}};
  _T_3323_im = _RAND_6136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6137 = {1{`RANDOM}};
  _T_3324_re = _RAND_6137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6138 = {1{`RANDOM}};
  _T_3324_im = _RAND_6138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6139 = {1{`RANDOM}};
  _T_3330_re = _RAND_6139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6140 = {1{`RANDOM}};
  _T_3330_im = _RAND_6140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6141 = {1{`RANDOM}};
  _T_3331_re = _RAND_6141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6142 = {1{`RANDOM}};
  _T_3331_im = _RAND_6142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6143 = {1{`RANDOM}};
  _T_3334_re = _RAND_6143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6144 = {1{`RANDOM}};
  _T_3334_im = _RAND_6144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6145 = {1{`RANDOM}};
  out1D1_re = _RAND_6145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6146 = {1{`RANDOM}};
  out1D1_im = _RAND_6146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6147 = {1{`RANDOM}};
  _T_3335_re = _RAND_6147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6148 = {1{`RANDOM}};
  _T_3335_im = _RAND_6148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6149 = {1{`RANDOM}};
  _T_3336_re = _RAND_6149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6150 = {1{`RANDOM}};
  _T_3336_im = _RAND_6150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 11'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    cntD1 <= cnt;
    cntD2 <= cntD1;
    out1_0_re <= io_dIn_re;
    out1_0_im <= io_dIn_im;
    out2_0_re <= io_dIn_re;
    out2_0_im <= io_dIn_im;
    _T_181_re <= out1_0_re;
    _T_181_im <= out1_0_im;
    _T_182_re <= _T_181_re;
    _T_182_im <= _T_181_im;
    _T_183_re <= _T_182_re;
    _T_183_im <= _T_182_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_325_re <= _T_324_re;
    _T_325_im <= _T_324_im;
    _T_326_re <= _T_325_re;
    _T_326_im <= _T_325_im;
    _T_327_re <= _T_326_re;
    _T_327_im <= _T_326_im;
    _T_328_re <= _T_327_re;
    _T_328_im <= _T_327_im;
    _T_329_re <= _T_328_re;
    _T_329_im <= _T_328_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_393_re <= _T_392_re;
    _T_393_im <= _T_392_im;
    _T_394_re <= _T_393_re;
    _T_394_im <= _T_393_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_402_re <= _T_401_re;
    _T_402_im <= _T_401_im;
    _T_403_re <= _T_402_re;
    _T_403_im <= _T_402_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_406_re <= _T_405_re;
    _T_406_im <= _T_405_im;
    _T_407_re <= _T_406_re;
    _T_407_im <= _T_406_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_409_re <= _T_408_re;
    _T_409_im <= _T_408_im;
    _T_410_re <= _T_409_re;
    _T_410_im <= _T_409_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_533_re <= _T_532_re;
    _T_533_im <= _T_532_im;
    _T_534_re <= _T_533_re;
    _T_534_im <= _T_533_im;
    _T_535_re <= _T_534_re;
    _T_535_im <= _T_534_im;
    _T_536_re <= _T_535_re;
    _T_536_im <= _T_535_im;
    _T_537_re <= _T_536_re;
    _T_537_im <= _T_536_im;
    _T_538_re <= _T_537_re;
    _T_538_im <= _T_537_im;
    _T_539_re <= _T_538_re;
    _T_539_im <= _T_538_im;
    _T_540_re <= _T_539_re;
    _T_540_im <= _T_539_im;
    _T_541_re <= _T_540_re;
    _T_541_im <= _T_540_im;
    _T_542_re <= _T_541_re;
    _T_542_im <= _T_541_im;
    _T_543_re <= _T_542_re;
    _T_543_im <= _T_542_im;
    _T_544_re <= _T_543_re;
    _T_544_im <= _T_543_im;
    _T_545_re <= _T_544_re;
    _T_545_im <= _T_544_im;
    _T_546_re <= _T_545_re;
    _T_546_im <= _T_545_im;
    _T_547_re <= _T_546_re;
    _T_547_im <= _T_546_im;
    _T_548_re <= _T_547_re;
    _T_548_im <= _T_547_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_663_re <= _T_662_re;
    _T_663_im <= _T_662_im;
    _T_664_re <= _T_663_re;
    _T_664_im <= _T_663_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_671_re <= _T_670_re;
    _T_671_im <= _T_670_im;
    _T_672_re <= _T_671_re;
    _T_672_im <= _T_671_im;
    _T_673_re <= _T_672_re;
    _T_673_im <= _T_672_im;
    _T_674_re <= _T_673_re;
    _T_674_im <= _T_673_im;
    _T_675_re <= _T_674_re;
    _T_675_im <= _T_674_im;
    _T_676_re <= _T_675_re;
    _T_676_im <= _T_675_im;
    _T_677_re <= _T_676_re;
    _T_677_im <= _T_676_im;
    _T_678_re <= _T_677_re;
    _T_678_im <= _T_677_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_728_re <= _T_727_re;
    _T_728_im <= _T_727_im;
    _T_729_re <= _T_728_re;
    _T_729_im <= _T_728_im;
    _T_730_re <= _T_729_re;
    _T_730_im <= _T_729_im;
    _T_731_re <= _T_730_re;
    _T_731_im <= _T_730_im;
    _T_732_re <= _T_731_re;
    _T_732_im <= _T_731_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_736_re <= _T_735_re;
    _T_736_im <= _T_735_im;
    _T_737_re <= _T_736_re;
    _T_737_im <= _T_736_im;
    _T_738_re <= _T_737_re;
    _T_738_im <= _T_737_im;
    _T_739_re <= _T_738_re;
    _T_739_im <= _T_738_im;
    _T_740_re <= _T_739_re;
    _T_740_im <= _T_739_im;
    _T_741_re <= _T_740_re;
    _T_741_im <= _T_740_im;
    _T_742_re <= _T_741_re;
    _T_742_im <= _T_741_im;
    _T_743_re <= _T_742_re;
    _T_743_im <= _T_742_im;
    _T_744_re <= _T_743_re;
    _T_744_im <= _T_743_im;
    _T_745_re <= _T_744_re;
    _T_745_im <= _T_744_im;
    _T_746_re <= _T_745_re;
    _T_746_im <= _T_745_im;
    _T_747_re <= _T_746_re;
    _T_747_im <= _T_746_im;
    _T_748_re <= _T_747_re;
    _T_748_im <= _T_747_im;
    _T_749_re <= _T_748_re;
    _T_749_im <= _T_748_im;
    _T_750_re <= _T_749_re;
    _T_750_im <= _T_749_im;
    _T_751_re <= _T_750_re;
    _T_751_im <= _T_750_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_796_re <= _T_795_re;
    _T_796_im <= _T_795_im;
    _T_797_re <= _T_796_re;
    _T_797_im <= _T_796_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_808_re <= _T_807_re;
    _T_808_im <= _T_807_im;
    _T_809_re <= _T_808_re;
    _T_809_im <= _T_808_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_811_re <= _T_810_re;
    _T_811_im <= _T_810_im;
    _T_812_re <= _T_811_re;
    _T_812_im <= _T_811_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_815_re <= _T_814_re;
    _T_815_im <= _T_814_im;
    _T_816_re <= _T_815_re;
    _T_816_im <= _T_815_im;
    _T_817_re <= _T_816_re;
    _T_817_im <= _T_816_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_829_re <= _T_828_re;
    _T_829_im <= _T_828_im;
    _T_830_re <= _T_829_re;
    _T_830_im <= _T_829_im;
    _T_831_re <= _T_830_re;
    _T_831_im <= _T_830_im;
    _T_832_re <= _T_831_re;
    _T_832_im <= _T_831_im;
    _T_833_re <= _T_832_re;
    _T_833_im <= _T_832_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_841_re <= _T_840_re;
    _T_841_im <= _T_840_im;
    _T_842_re <= _T_841_re;
    _T_842_im <= _T_841_im;
    _T_843_re <= _T_842_re;
    _T_843_im <= _T_842_im;
    _T_844_re <= _T_843_re;
    _T_844_im <= _T_843_im;
    _T_845_re <= _T_844_re;
    _T_845_im <= _T_844_im;
    _T_846_re <= _T_845_re;
    _T_846_im <= _T_845_im;
    _T_847_re <= _T_846_re;
    _T_847_im <= _T_846_im;
    _T_848_re <= _T_847_re;
    _T_848_im <= _T_847_im;
    _T_849_re <= _T_848_re;
    _T_849_im <= _T_848_im;
    _T_850_re <= _T_849_re;
    _T_850_im <= _T_849_im;
    _T_851_re <= _T_850_re;
    _T_851_im <= _T_850_im;
    _T_852_re <= _T_851_re;
    _T_852_im <= _T_851_im;
    _T_853_re <= _T_852_re;
    _T_853_im <= _T_852_im;
    _T_854_re <= _T_853_re;
    _T_854_im <= _T_853_im;
    _T_855_re <= _T_854_re;
    _T_855_im <= _T_854_im;
    _T_856_re <= _T_855_re;
    _T_856_im <= _T_855_im;
    _T_857_re <= _T_856_re;
    _T_857_im <= _T_856_im;
    _T_858_re <= _T_857_re;
    _T_858_im <= _T_857_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_865_re <= _T_864_re;
    _T_865_im <= _T_864_im;
    _T_866_re <= _T_865_re;
    _T_866_im <= _T_865_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_881_re <= _T_880_re;
    _T_881_im <= _T_880_im;
    _T_882_re <= _T_881_re;
    _T_882_im <= _T_881_im;
    _T_883_re <= _T_882_re;
    _T_883_im <= _T_882_im;
    _T_884_re <= _T_883_re;
    _T_884_im <= _T_883_im;
    _T_885_re <= _T_884_re;
    _T_885_im <= _T_884_im;
    _T_886_re <= _T_885_re;
    _T_886_im <= _T_885_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_890_re <= _T_889_re;
    _T_890_im <= _T_889_im;
    _T_891_re <= _T_890_re;
    _T_891_im <= _T_890_im;
    _T_892_re <= _T_891_re;
    _T_892_im <= _T_891_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_898_re <= _T_897_re;
    _T_898_im <= _T_897_im;
    _T_899_re <= _T_898_re;
    _T_899_im <= _T_898_im;
    _T_900_re <= _T_899_re;
    _T_900_im <= _T_899_im;
    _T_901_re <= _T_900_re;
    _T_901_im <= _T_900_im;
    _T_902_re <= _T_901_re;
    _T_902_im <= _T_901_im;
    _T_903_re <= _T_902_re;
    _T_903_im <= _T_902_im;
    _T_904_re <= _T_903_re;
    _T_904_im <= _T_903_im;
    _T_905_re <= _T_904_re;
    _T_905_im <= _T_904_im;
    _T_906_re <= _T_905_re;
    _T_906_im <= _T_905_im;
    _T_907_re <= _T_906_re;
    _T_907_im <= _T_906_im;
    _T_908_re <= _T_907_re;
    _T_908_im <= _T_907_im;
    _T_909_re <= _T_908_re;
    _T_909_im <= _T_908_im;
    _T_910_re <= _T_909_re;
    _T_910_im <= _T_909_im;
    _T_911_re <= _T_910_re;
    _T_911_im <= _T_910_im;
    _T_912_re <= _T_911_re;
    _T_912_im <= _T_911_im;
    _T_913_re <= _T_912_re;
    _T_913_im <= _T_912_im;
    _T_914_re <= _T_913_re;
    _T_914_im <= _T_913_im;
    _T_915_re <= _T_914_re;
    _T_915_im <= _T_914_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_922_re <= _T_921_re;
    _T_922_im <= _T_921_im;
    _T_923_re <= _T_922_re;
    _T_923_im <= _T_922_im;
    _T_924_re <= _T_923_re;
    _T_924_im <= _T_923_im;
    _T_925_re <= _T_924_re;
    _T_925_im <= _T_924_im;
    _T_926_re <= _T_925_re;
    _T_926_im <= _T_925_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_928_re <= _T_927_re;
    _T_928_im <= _T_927_im;
    _T_929_re <= _T_928_re;
    _T_929_im <= _T_928_im;
    _T_930_re <= _T_929_re;
    _T_930_im <= _T_929_im;
    _T_931_re <= _T_930_re;
    _T_931_im <= _T_930_im;
    _T_932_re <= _T_931_re;
    _T_932_im <= _T_931_im;
    _T_933_re <= _T_932_re;
    _T_933_im <= _T_932_im;
    _T_934_re <= _T_933_re;
    _T_934_im <= _T_933_im;
    _T_935_re <= _T_934_re;
    _T_935_im <= _T_934_im;
    _T_936_re <= _T_935_re;
    _T_936_im <= _T_935_im;
    _T_937_re <= _T_936_re;
    _T_937_im <= _T_936_im;
    _T_938_re <= _T_937_re;
    _T_938_im <= _T_937_im;
    _T_939_re <= _T_938_re;
    _T_939_im <= _T_938_im;
    _T_940_re <= _T_939_re;
    _T_940_im <= _T_939_im;
    _T_941_re <= _T_940_re;
    _T_941_im <= _T_940_im;
    _T_942_re <= _T_941_re;
    _T_942_im <= _T_941_im;
    _T_943_re <= _T_942_re;
    _T_943_im <= _T_942_im;
    _T_944_re <= _T_943_re;
    _T_944_im <= _T_943_im;
    _T_945_re <= _T_944_re;
    _T_945_im <= _T_944_im;
    _T_946_re <= _T_945_re;
    _T_946_im <= _T_945_im;
    _T_947_re <= _T_946_re;
    _T_947_im <= _T_946_im;
    _T_948_re <= _T_947_re;
    _T_948_im <= _T_947_im;
    _T_949_re <= _T_948_re;
    _T_949_im <= _T_948_im;
    _T_950_re <= _T_949_re;
    _T_950_im <= _T_949_im;
    _T_951_re <= _T_950_re;
    _T_951_im <= _T_950_im;
    _T_952_re <= _T_951_re;
    _T_952_im <= _T_951_im;
    _T_953_re <= _T_952_re;
    _T_953_im <= _T_952_im;
    _T_954_re <= _T_953_re;
    _T_954_im <= _T_953_im;
    _T_955_re <= _T_954_re;
    _T_955_im <= _T_954_im;
    _T_956_re <= _T_955_re;
    _T_956_im <= _T_955_im;
    _T_957_re <= _T_956_re;
    _T_957_im <= _T_956_im;
    _T_958_re <= _T_957_re;
    _T_958_im <= _T_957_im;
    _T_959_re <= _T_958_re;
    _T_959_im <= _T_958_im;
    _T_960_re <= _T_959_re;
    _T_960_im <= _T_959_im;
    _T_961_re <= _T_960_re;
    _T_961_im <= _T_960_im;
    _T_962_re <= _T_961_re;
    _T_962_im <= _T_961_im;
    _T_963_re <= _T_962_re;
    _T_963_im <= _T_962_im;
    _T_964_re <= _T_963_re;
    _T_964_im <= _T_963_im;
    _T_965_re <= _T_964_re;
    _T_965_im <= _T_964_im;
    _T_966_re <= _T_965_re;
    _T_966_im <= _T_965_im;
    _T_967_re <= _T_966_re;
    _T_967_im <= _T_966_im;
    _T_968_re <= _T_967_re;
    _T_968_im <= _T_967_im;
    _T_969_re <= _T_968_re;
    _T_969_im <= _T_968_im;
    _T_970_re <= _T_969_re;
    _T_970_im <= _T_969_im;
    _T_971_re <= _T_970_re;
    _T_971_im <= _T_970_im;
    _T_972_re <= _T_971_re;
    _T_972_im <= _T_971_im;
    _T_973_re <= _T_972_re;
    _T_973_im <= _T_972_im;
    _T_974_re <= _T_973_re;
    _T_974_im <= _T_973_im;
    _T_975_re <= _T_974_re;
    _T_975_im <= _T_974_im;
    _T_976_re <= _T_975_re;
    _T_976_im <= _T_975_im;
    _T_977_re <= _T_976_re;
    _T_977_im <= _T_976_im;
    _T_978_re <= _T_977_re;
    _T_978_im <= _T_977_im;
    _T_979_re <= _T_978_re;
    _T_979_im <= _T_978_im;
    _T_980_re <= _T_979_re;
    _T_980_im <= _T_979_im;
    _T_981_re <= _T_980_re;
    _T_981_im <= _T_980_im;
    _T_982_re <= _T_981_re;
    _T_982_im <= _T_981_im;
    _T_983_re <= _T_982_re;
    _T_983_im <= _T_982_im;
    _T_984_re <= _T_983_re;
    _T_984_im <= _T_983_im;
    _T_985_re <= _T_984_re;
    _T_985_im <= _T_984_im;
    _T_986_re <= _T_985_re;
    _T_986_im <= _T_985_im;
    _T_987_re <= _T_986_re;
    _T_987_im <= _T_986_im;
    _T_988_re <= _T_987_re;
    _T_988_im <= _T_987_im;
    _T_989_re <= _T_988_re;
    _T_989_im <= _T_988_im;
    _T_990_re <= _T_989_re;
    _T_990_im <= _T_989_im;
    _T_991_re <= _T_990_re;
    _T_991_im <= _T_990_im;
    _T_992_re <= _T_991_re;
    _T_992_im <= _T_991_im;
    _T_993_re <= _T_992_re;
    _T_993_im <= _T_992_im;
    _T_994_re <= _T_993_re;
    _T_994_im <= _T_993_im;
    _T_995_re <= _T_994_re;
    _T_995_im <= _T_994_im;
    _T_996_re <= _T_995_re;
    _T_996_im <= _T_995_im;
    _T_997_re <= _T_996_re;
    _T_997_im <= _T_996_im;
    _T_998_re <= _T_997_re;
    _T_998_im <= _T_997_im;
    _T_999_re <= _T_998_re;
    _T_999_im <= _T_998_im;
    _T_1000_re <= _T_999_re;
    _T_1000_im <= _T_999_im;
    _T_1001_re <= _T_1000_re;
    _T_1001_im <= _T_1000_im;
    _T_1002_re <= _T_1001_re;
    _T_1002_im <= _T_1001_im;
    _T_1003_re <= _T_1002_re;
    _T_1003_im <= _T_1002_im;
    _T_1004_re <= _T_1003_re;
    _T_1004_im <= _T_1003_im;
    _T_1005_re <= _T_1004_re;
    _T_1005_im <= _T_1004_im;
    _T_1006_re <= _T_1005_re;
    _T_1006_im <= _T_1005_im;
    _T_1007_re <= _T_1006_re;
    _T_1007_im <= _T_1006_im;
    _T_1008_re <= _T_1007_re;
    _T_1008_im <= _T_1007_im;
    _T_1009_re <= _T_1008_re;
    _T_1009_im <= _T_1008_im;
    _T_1010_re <= _T_1009_re;
    _T_1010_im <= _T_1009_im;
    _T_1011_re <= _T_1010_re;
    _T_1011_im <= _T_1010_im;
    _T_1012_re <= _T_1011_re;
    _T_1012_im <= _T_1011_im;
    _T_1013_re <= _T_1012_re;
    _T_1013_im <= _T_1012_im;
    _T_1014_re <= _T_1013_re;
    _T_1014_im <= _T_1013_im;
    _T_1015_re <= _T_1014_re;
    _T_1015_im <= _T_1014_im;
    _T_1016_re <= _T_1015_re;
    _T_1016_im <= _T_1015_im;
    _T_1017_re <= _T_1016_re;
    _T_1017_im <= _T_1016_im;
    _T_1018_re <= _T_1017_re;
    _T_1018_im <= _T_1017_im;
    _T_1019_re <= _T_1018_re;
    _T_1019_im <= _T_1018_im;
    _T_1020_re <= _T_1019_re;
    _T_1020_im <= _T_1019_im;
    _T_1021_re <= _T_1020_re;
    _T_1021_im <= _T_1020_im;
    _T_1022_re <= _T_1021_re;
    _T_1022_im <= _T_1021_im;
    _T_1023_re <= _T_1022_re;
    _T_1023_im <= _T_1022_im;
    _T_1024_re <= _T_1023_re;
    _T_1024_im <= _T_1023_im;
    _T_1025_re <= _T_1024_re;
    _T_1025_im <= _T_1024_im;
    _T_1026_re <= _T_1025_re;
    _T_1026_im <= _T_1025_im;
    _T_1027_re <= _T_1026_re;
    _T_1027_im <= _T_1026_im;
    _T_1028_re <= _T_1027_re;
    _T_1028_im <= _T_1027_im;
    _T_1029_re <= _T_1028_re;
    _T_1029_im <= _T_1028_im;
    _T_1030_re <= _T_1029_re;
    _T_1030_im <= _T_1029_im;
    _T_1031_re <= _T_1030_re;
    _T_1031_im <= _T_1030_im;
    _T_1032_re <= _T_1031_re;
    _T_1032_im <= _T_1031_im;
    _T_1033_re <= _T_1032_re;
    _T_1033_im <= _T_1032_im;
    _T_1034_re <= _T_1033_re;
    _T_1034_im <= _T_1033_im;
    _T_1035_re <= _T_1034_re;
    _T_1035_im <= _T_1034_im;
    _T_1036_re <= _T_1035_re;
    _T_1036_im <= _T_1035_im;
    _T_1037_re <= _T_1036_re;
    _T_1037_im <= _T_1036_im;
    _T_1038_re <= _T_1037_re;
    _T_1038_im <= _T_1037_im;
    _T_1039_re <= _T_1038_re;
    _T_1039_im <= _T_1038_im;
    _T_1040_re <= _T_1039_re;
    _T_1040_im <= _T_1039_im;
    _T_1041_re <= _T_1040_re;
    _T_1041_im <= _T_1040_im;
    _T_1042_re <= _T_1041_re;
    _T_1042_im <= _T_1041_im;
    _T_1043_re <= _T_1042_re;
    _T_1043_im <= _T_1042_im;
    _T_1044_re <= _T_1043_re;
    _T_1044_im <= _T_1043_im;
    _T_1045_re <= _T_1044_re;
    _T_1045_im <= _T_1044_im;
    _T_1046_re <= _T_1045_re;
    _T_1046_im <= _T_1045_im;
    _T_1047_re <= _T_1046_re;
    _T_1047_im <= _T_1046_im;
    _T_1048_re <= _T_1047_re;
    _T_1048_im <= _T_1047_im;
    _T_1049_re <= _T_1048_re;
    _T_1049_im <= _T_1048_im;
    _T_1050_re <= _T_1049_re;
    _T_1050_im <= _T_1049_im;
    _T_1051_re <= _T_1050_re;
    _T_1051_im <= _T_1050_im;
    _T_1052_re <= _T_1051_re;
    _T_1052_im <= _T_1051_im;
    _T_1053_re <= _T_1052_re;
    _T_1053_im <= _T_1052_im;
    _T_1054_re <= _T_1053_re;
    _T_1054_im <= _T_1053_im;
    _T_1055_re <= _T_1054_re;
    _T_1055_im <= _T_1054_im;
    _T_1056_re <= _T_1055_re;
    _T_1056_im <= _T_1055_im;
    _T_1057_re <= _T_1056_re;
    _T_1057_im <= _T_1056_im;
    _T_1058_re <= _T_1057_re;
    _T_1058_im <= _T_1057_im;
    _T_1059_re <= _T_1058_re;
    _T_1059_im <= _T_1058_im;
    _T_1060_re <= _T_1059_re;
    _T_1060_im <= _T_1059_im;
    _T_1061_re <= _T_1060_re;
    _T_1061_im <= _T_1060_im;
    _T_1062_re <= _T_1061_re;
    _T_1062_im <= _T_1061_im;
    _T_1063_re <= _T_1062_re;
    _T_1063_im <= _T_1062_im;
    _T_1064_re <= _T_1063_re;
    _T_1064_im <= _T_1063_im;
    _T_1065_re <= _T_1064_re;
    _T_1065_im <= _T_1064_im;
    _T_1066_re <= _T_1065_re;
    _T_1066_im <= _T_1065_im;
    _T_1067_re <= _T_1066_re;
    _T_1067_im <= _T_1066_im;
    _T_1068_re <= _T_1067_re;
    _T_1068_im <= _T_1067_im;
    _T_1069_re <= _T_1068_re;
    _T_1069_im <= _T_1068_im;
    _T_1070_re <= _T_1069_re;
    _T_1070_im <= _T_1069_im;
    _T_1071_re <= _T_1070_re;
    _T_1071_im <= _T_1070_im;
    _T_1072_re <= _T_1071_re;
    _T_1072_im <= _T_1071_im;
    _T_1073_re <= _T_1072_re;
    _T_1073_im <= _T_1072_im;
    _T_1074_re <= _T_1073_re;
    _T_1074_im <= _T_1073_im;
    _T_1075_re <= _T_1074_re;
    _T_1075_im <= _T_1074_im;
    _T_1076_re <= _T_1075_re;
    _T_1076_im <= _T_1075_im;
    _T_1077_re <= _T_1076_re;
    _T_1077_im <= _T_1076_im;
    _T_1078_re <= _T_1077_re;
    _T_1078_im <= _T_1077_im;
    _T_1079_re <= _T_1078_re;
    _T_1079_im <= _T_1078_im;
    _T_1080_re <= _T_1079_re;
    _T_1080_im <= _T_1079_im;
    _T_1081_re <= _T_1080_re;
    _T_1081_im <= _T_1080_im;
    _T_1082_re <= _T_1081_re;
    _T_1082_im <= _T_1081_im;
    _T_1083_re <= _T_1082_re;
    _T_1083_im <= _T_1082_im;
    _T_1084_re <= _T_1083_re;
    _T_1084_im <= _T_1083_im;
    _T_1085_re <= _T_1084_re;
    _T_1085_im <= _T_1084_im;
    _T_1086_re <= _T_1085_re;
    _T_1086_im <= _T_1085_im;
    _T_1087_re <= _T_1086_re;
    _T_1087_im <= _T_1086_im;
    _T_1088_re <= _T_1087_re;
    _T_1088_im <= _T_1087_im;
    _T_1089_re <= _T_1088_re;
    _T_1089_im <= _T_1088_im;
    _T_1090_re <= _T_1089_re;
    _T_1090_im <= _T_1089_im;
    _T_1091_re <= _T_1090_re;
    _T_1091_im <= _T_1090_im;
    _T_1092_re <= _T_1091_re;
    _T_1092_im <= _T_1091_im;
    _T_1093_re <= _T_1092_re;
    _T_1093_im <= _T_1092_im;
    _T_1094_re <= _T_1093_re;
    _T_1094_im <= _T_1093_im;
    _T_1095_re <= _T_1094_re;
    _T_1095_im <= _T_1094_im;
    _T_1096_re <= _T_1095_re;
    _T_1096_im <= _T_1095_im;
    _T_1097_re <= _T_1096_re;
    _T_1097_im <= _T_1096_im;
    _T_1098_re <= _T_1097_re;
    _T_1098_im <= _T_1097_im;
    _T_1099_re <= _T_1098_re;
    _T_1099_im <= _T_1098_im;
    _T_1100_re <= _T_1099_re;
    _T_1100_im <= _T_1099_im;
    _T_1101_re <= _T_1100_re;
    _T_1101_im <= _T_1100_im;
    _T_1102_re <= _T_1101_re;
    _T_1102_im <= _T_1101_im;
    _T_1103_re <= _T_1102_re;
    _T_1103_im <= _T_1102_im;
    _T_1104_re <= _T_1103_re;
    _T_1104_im <= _T_1103_im;
    _T_1105_re <= _T_1104_re;
    _T_1105_im <= _T_1104_im;
    _T_1106_re <= _T_1105_re;
    _T_1106_im <= _T_1105_im;
    _T_1107_re <= _T_1106_re;
    _T_1107_im <= _T_1106_im;
    _T_1108_re <= _T_1107_re;
    _T_1108_im <= _T_1107_im;
    _T_1109_re <= _T_1108_re;
    _T_1109_im <= _T_1108_im;
    _T_1110_re <= _T_1109_re;
    _T_1110_im <= _T_1109_im;
    _T_1111_re <= _T_1110_re;
    _T_1111_im <= _T_1110_im;
    _T_1112_re <= _T_1111_re;
    _T_1112_im <= _T_1111_im;
    _T_1113_re <= _T_1112_re;
    _T_1113_im <= _T_1112_im;
    _T_1114_re <= _T_1113_re;
    _T_1114_im <= _T_1113_im;
    _T_1115_re <= _T_1114_re;
    _T_1115_im <= _T_1114_im;
    _T_1116_re <= _T_1115_re;
    _T_1116_im <= _T_1115_im;
    _T_1117_re <= _T_1116_re;
    _T_1117_im <= _T_1116_im;
    _T_1118_re <= _T_1117_re;
    _T_1118_im <= _T_1117_im;
    _T_1119_re <= _T_1118_re;
    _T_1119_im <= _T_1118_im;
    _T_1120_re <= _T_1119_re;
    _T_1120_im <= _T_1119_im;
    _T_1121_re <= _T_1120_re;
    _T_1121_im <= _T_1120_im;
    _T_1122_re <= _T_1121_re;
    _T_1122_im <= _T_1121_im;
    _T_1123_re <= _T_1122_re;
    _T_1123_im <= _T_1122_im;
    _T_1124_re <= _T_1123_re;
    _T_1124_im <= _T_1123_im;
    _T_1125_re <= _T_1124_re;
    _T_1125_im <= _T_1124_im;
    _T_1126_re <= _T_1125_re;
    _T_1126_im <= _T_1125_im;
    _T_1127_re <= _T_1126_re;
    _T_1127_im <= _T_1126_im;
    _T_1128_re <= _T_1127_re;
    _T_1128_im <= _T_1127_im;
    _T_1129_re <= _T_1128_re;
    _T_1129_im <= _T_1128_im;
    _T_1130_re <= _T_1129_re;
    _T_1130_im <= _T_1129_im;
    _T_1131_re <= _T_1130_re;
    _T_1131_im <= _T_1130_im;
    _T_1132_re <= _T_1131_re;
    _T_1132_im <= _T_1131_im;
    _T_1133_re <= _T_1132_re;
    _T_1133_im <= _T_1132_im;
    _T_1134_re <= _T_1133_re;
    _T_1134_im <= _T_1133_im;
    _T_1135_re <= _T_1134_re;
    _T_1135_im <= _T_1134_im;
    _T_1136_re <= _T_1135_re;
    _T_1136_im <= _T_1135_im;
    _T_1137_re <= _T_1136_re;
    _T_1137_im <= _T_1136_im;
    _T_1138_re <= _T_1137_re;
    _T_1138_im <= _T_1137_im;
    _T_1139_re <= _T_1138_re;
    _T_1139_im <= _T_1138_im;
    _T_1140_re <= _T_1139_re;
    _T_1140_im <= _T_1139_im;
    _T_1141_re <= _T_1140_re;
    _T_1141_im <= _T_1140_im;
    _T_1142_re <= _T_1141_re;
    _T_1142_im <= _T_1141_im;
    _T_1143_re <= _T_1142_re;
    _T_1143_im <= _T_1142_im;
    _T_1144_re <= _T_1143_re;
    _T_1144_im <= _T_1143_im;
    _T_1145_re <= _T_1144_re;
    _T_1145_im <= _T_1144_im;
    _T_1146_re <= _T_1145_re;
    _T_1146_im <= _T_1145_im;
    _T_1147_re <= _T_1146_re;
    _T_1147_im <= _T_1146_im;
    _T_1148_re <= _T_1147_re;
    _T_1148_im <= _T_1147_im;
    _T_1149_re <= _T_1148_re;
    _T_1149_im <= _T_1148_im;
    _T_1150_re <= _T_1149_re;
    _T_1150_im <= _T_1149_im;
    _T_1151_re <= _T_1150_re;
    _T_1151_im <= _T_1150_im;
    _T_1152_re <= _T_1151_re;
    _T_1152_im <= _T_1151_im;
    _T_1153_re <= _T_1152_re;
    _T_1153_im <= _T_1152_im;
    _T_1154_re <= _T_1153_re;
    _T_1154_im <= _T_1153_im;
    _T_1155_re <= _T_1154_re;
    _T_1155_im <= _T_1154_im;
    _T_1156_re <= _T_1155_re;
    _T_1156_im <= _T_1155_im;
    _T_1157_re <= _T_1156_re;
    _T_1157_im <= _T_1156_im;
    _T_1158_re <= _T_1157_re;
    _T_1158_im <= _T_1157_im;
    _T_1159_re <= _T_1158_re;
    _T_1159_im <= _T_1158_im;
    _T_1160_re <= _T_1159_re;
    _T_1160_im <= _T_1159_im;
    _T_1161_re <= _T_1160_re;
    _T_1161_im <= _T_1160_im;
    _T_1162_re <= _T_1161_re;
    _T_1162_im <= _T_1161_im;
    _T_1163_re <= _T_1162_re;
    _T_1163_im <= _T_1162_im;
    _T_1164_re <= _T_1163_re;
    _T_1164_im <= _T_1163_im;
    _T_1165_re <= _T_1164_re;
    _T_1165_im <= _T_1164_im;
    _T_1166_re <= _T_1165_re;
    _T_1166_im <= _T_1165_im;
    _T_1167_re <= _T_1166_re;
    _T_1167_im <= _T_1166_im;
    _T_1168_re <= _T_1167_re;
    _T_1168_im <= _T_1167_im;
    _T_1169_re <= _T_1168_re;
    _T_1169_im <= _T_1168_im;
    _T_1170_re <= _T_1169_re;
    _T_1170_im <= _T_1169_im;
    _T_1171_re <= _T_1170_re;
    _T_1171_im <= _T_1170_im;
    _T_1172_re <= _T_1171_re;
    _T_1172_im <= _T_1171_im;
    _T_1173_re <= _T_1172_re;
    _T_1173_im <= _T_1172_im;
    _T_1174_re <= _T_1173_re;
    _T_1174_im <= _T_1173_im;
    _T_1175_re <= _T_1174_re;
    _T_1175_im <= _T_1174_im;
    _T_1176_re <= _T_1175_re;
    _T_1176_im <= _T_1175_im;
    _T_1177_re <= _T_1176_re;
    _T_1177_im <= _T_1176_im;
    _T_1178_re <= _T_1177_re;
    _T_1178_im <= _T_1177_im;
    _T_1179_re <= _T_1178_re;
    _T_1179_im <= _T_1178_im;
    _T_1180_re <= _T_1179_re;
    _T_1180_im <= _T_1179_im;
    _T_1181_re <= _T_1180_re;
    _T_1181_im <= _T_1180_im;
    _T_1182_re <= _T_1181_re;
    _T_1182_im <= _T_1181_im;
    _T_1183_re <= _T_1182_re;
    _T_1183_im <= _T_1182_im;
    _T_1184_re <= _T_1183_re;
    _T_1184_im <= _T_1183_im;
    _T_1185_re <= _T_1184_re;
    _T_1185_im <= _T_1184_im;
    _T_1186_re <= _T_1185_re;
    _T_1186_im <= _T_1185_im;
    _T_1187_re <= _T_1186_re;
    _T_1187_im <= _T_1186_im;
    _T_1188_re <= _T_1187_re;
    _T_1188_im <= _T_1187_im;
    _T_1189_re <= _T_1188_re;
    _T_1189_im <= _T_1188_im;
    _T_1190_re <= _T_1189_re;
    _T_1190_im <= _T_1189_im;
    _T_1191_re <= _T_1190_re;
    _T_1191_im <= _T_1190_im;
    _T_1192_re <= _T_1191_re;
    _T_1192_im <= _T_1191_im;
    _T_1193_re <= _T_1192_re;
    _T_1193_im <= _T_1192_im;
    _T_1194_re <= _T_1193_re;
    _T_1194_im <= _T_1193_im;
    _T_1195_re <= _T_1194_re;
    _T_1195_im <= _T_1194_im;
    _T_1196_re <= _T_1195_re;
    _T_1196_im <= _T_1195_im;
    _T_1197_re <= _T_1196_re;
    _T_1197_im <= _T_1196_im;
    _T_1198_re <= _T_1197_re;
    _T_1198_im <= _T_1197_im;
    _T_1199_re <= _T_1198_re;
    _T_1199_im <= _T_1198_im;
    _T_1200_re <= _T_1199_re;
    _T_1200_im <= _T_1199_im;
    _T_1201_re <= _T_1200_re;
    _T_1201_im <= _T_1200_im;
    _T_1202_re <= _T_1201_re;
    _T_1202_im <= _T_1201_im;
    _T_1203_re <= _T_1202_re;
    _T_1203_im <= _T_1202_im;
    _T_1204_re <= _T_1203_re;
    _T_1204_im <= _T_1203_im;
    _T_1207_re <= Butterfly_io_out2_re;
    _T_1207_im <= Butterfly_io_out2_im;
    _T_1208_re <= _T_1207_re;
    _T_1208_im <= _T_1207_im;
    _T_1209_re <= _T_1208_re;
    _T_1209_im <= _T_1208_im;
    _T_1210_re <= _T_1209_re;
    _T_1210_im <= _T_1209_im;
    _T_1211_re <= _T_1210_re;
    _T_1211_im <= _T_1210_im;
    _T_1212_re <= _T_1211_re;
    _T_1212_im <= _T_1211_im;
    _T_1213_re <= _T_1212_re;
    _T_1213_im <= _T_1212_im;
    _T_1214_re <= _T_1213_re;
    _T_1214_im <= _T_1213_im;
    _T_1215_re <= _T_1214_re;
    _T_1215_im <= _T_1214_im;
    _T_1216_re <= _T_1215_re;
    _T_1216_im <= _T_1215_im;
    _T_1217_re <= _T_1216_re;
    _T_1217_im <= _T_1216_im;
    _T_1218_re <= _T_1217_re;
    _T_1218_im <= _T_1217_im;
    _T_1219_re <= _T_1218_re;
    _T_1219_im <= _T_1218_im;
    _T_1220_re <= _T_1219_re;
    _T_1220_im <= _T_1219_im;
    _T_1221_re <= _T_1220_re;
    _T_1221_im <= _T_1220_im;
    _T_1222_re <= _T_1221_re;
    _T_1222_im <= _T_1221_im;
    _T_1223_re <= _T_1222_re;
    _T_1223_im <= _T_1222_im;
    _T_1224_re <= _T_1223_re;
    _T_1224_im <= _T_1223_im;
    _T_1225_re <= _T_1224_re;
    _T_1225_im <= _T_1224_im;
    _T_1226_re <= _T_1225_re;
    _T_1226_im <= _T_1225_im;
    _T_1227_re <= _T_1226_re;
    _T_1227_im <= _T_1226_im;
    _T_1228_re <= _T_1227_re;
    _T_1228_im <= _T_1227_im;
    _T_1229_re <= _T_1228_re;
    _T_1229_im <= _T_1228_im;
    _T_1230_re <= _T_1229_re;
    _T_1230_im <= _T_1229_im;
    _T_1231_re <= _T_1230_re;
    _T_1231_im <= _T_1230_im;
    _T_1232_re <= _T_1231_re;
    _T_1232_im <= _T_1231_im;
    _T_1233_re <= _T_1232_re;
    _T_1233_im <= _T_1232_im;
    _T_1234_re <= _T_1233_re;
    _T_1234_im <= _T_1233_im;
    _T_1235_re <= _T_1234_re;
    _T_1235_im <= _T_1234_im;
    _T_1236_re <= _T_1235_re;
    _T_1236_im <= _T_1235_im;
    _T_1237_re <= _T_1236_re;
    _T_1237_im <= _T_1236_im;
    _T_1238_re <= _T_1237_re;
    _T_1238_im <= _T_1237_im;
    _T_1239_re <= _T_1238_re;
    _T_1239_im <= _T_1238_im;
    _T_1240_re <= _T_1239_re;
    _T_1240_im <= _T_1239_im;
    _T_1241_re <= _T_1240_re;
    _T_1241_im <= _T_1240_im;
    _T_1242_re <= _T_1241_re;
    _T_1242_im <= _T_1241_im;
    _T_1243_re <= _T_1242_re;
    _T_1243_im <= _T_1242_im;
    _T_1244_re <= _T_1243_re;
    _T_1244_im <= _T_1243_im;
    _T_1245_re <= _T_1244_re;
    _T_1245_im <= _T_1244_im;
    _T_1246_re <= _T_1245_re;
    _T_1246_im <= _T_1245_im;
    _T_1247_re <= _T_1246_re;
    _T_1247_im <= _T_1246_im;
    _T_1248_re <= _T_1247_re;
    _T_1248_im <= _T_1247_im;
    _T_1249_re <= _T_1248_re;
    _T_1249_im <= _T_1248_im;
    _T_1250_re <= _T_1249_re;
    _T_1250_im <= _T_1249_im;
    _T_1251_re <= _T_1250_re;
    _T_1251_im <= _T_1250_im;
    _T_1252_re <= _T_1251_re;
    _T_1252_im <= _T_1251_im;
    _T_1253_re <= _T_1252_re;
    _T_1253_im <= _T_1252_im;
    _T_1254_re <= _T_1253_re;
    _T_1254_im <= _T_1253_im;
    _T_1255_re <= _T_1254_re;
    _T_1255_im <= _T_1254_im;
    _T_1256_re <= _T_1255_re;
    _T_1256_im <= _T_1255_im;
    _T_1257_re <= _T_1256_re;
    _T_1257_im <= _T_1256_im;
    _T_1258_re <= _T_1257_re;
    _T_1258_im <= _T_1257_im;
    _T_1259_re <= _T_1258_re;
    _T_1259_im <= _T_1258_im;
    _T_1260_re <= _T_1259_re;
    _T_1260_im <= _T_1259_im;
    _T_1261_re <= _T_1260_re;
    _T_1261_im <= _T_1260_im;
    _T_1262_re <= _T_1261_re;
    _T_1262_im <= _T_1261_im;
    _T_1263_re <= _T_1262_re;
    _T_1263_im <= _T_1262_im;
    _T_1264_re <= _T_1263_re;
    _T_1264_im <= _T_1263_im;
    _T_1265_re <= _T_1264_re;
    _T_1265_im <= _T_1264_im;
    _T_1266_re <= _T_1265_re;
    _T_1266_im <= _T_1265_im;
    _T_1267_re <= _T_1266_re;
    _T_1267_im <= _T_1266_im;
    _T_1268_re <= _T_1267_re;
    _T_1268_im <= _T_1267_im;
    _T_1269_re <= _T_1268_re;
    _T_1269_im <= _T_1268_im;
    _T_1270_re <= _T_1269_re;
    _T_1270_im <= _T_1269_im;
    _T_1271_re <= _T_1270_re;
    _T_1271_im <= _T_1270_im;
    _T_1272_re <= _T_1271_re;
    _T_1272_im <= _T_1271_im;
    _T_1273_re <= _T_1272_re;
    _T_1273_im <= _T_1272_im;
    _T_1274_re <= _T_1273_re;
    _T_1274_im <= _T_1273_im;
    _T_1275_re <= _T_1274_re;
    _T_1275_im <= _T_1274_im;
    _T_1276_re <= _T_1275_re;
    _T_1276_im <= _T_1275_im;
    _T_1277_re <= _T_1276_re;
    _T_1277_im <= _T_1276_im;
    _T_1278_re <= _T_1277_re;
    _T_1278_im <= _T_1277_im;
    _T_1279_re <= _T_1278_re;
    _T_1279_im <= _T_1278_im;
    _T_1280_re <= _T_1279_re;
    _T_1280_im <= _T_1279_im;
    _T_1281_re <= _T_1280_re;
    _T_1281_im <= _T_1280_im;
    _T_1282_re <= _T_1281_re;
    _T_1282_im <= _T_1281_im;
    _T_1283_re <= _T_1282_re;
    _T_1283_im <= _T_1282_im;
    _T_1284_re <= _T_1283_re;
    _T_1284_im <= _T_1283_im;
    _T_1285_re <= _T_1284_re;
    _T_1285_im <= _T_1284_im;
    _T_1286_re <= _T_1285_re;
    _T_1286_im <= _T_1285_im;
    _T_1287_re <= _T_1286_re;
    _T_1287_im <= _T_1286_im;
    _T_1288_re <= _T_1287_re;
    _T_1288_im <= _T_1287_im;
    _T_1289_re <= _T_1288_re;
    _T_1289_im <= _T_1288_im;
    _T_1290_re <= _T_1289_re;
    _T_1290_im <= _T_1289_im;
    _T_1291_re <= _T_1290_re;
    _T_1291_im <= _T_1290_im;
    _T_1292_re <= _T_1291_re;
    _T_1292_im <= _T_1291_im;
    _T_1293_re <= _T_1292_re;
    _T_1293_im <= _T_1292_im;
    _T_1294_re <= _T_1293_re;
    _T_1294_im <= _T_1293_im;
    _T_1295_re <= _T_1294_re;
    _T_1295_im <= _T_1294_im;
    _T_1296_re <= _T_1295_re;
    _T_1296_im <= _T_1295_im;
    _T_1297_re <= _T_1296_re;
    _T_1297_im <= _T_1296_im;
    _T_1298_re <= _T_1297_re;
    _T_1298_im <= _T_1297_im;
    _T_1299_re <= _T_1298_re;
    _T_1299_im <= _T_1298_im;
    _T_1300_re <= _T_1299_re;
    _T_1300_im <= _T_1299_im;
    _T_1301_re <= _T_1300_re;
    _T_1301_im <= _T_1300_im;
    _T_1302_re <= _T_1301_re;
    _T_1302_im <= _T_1301_im;
    _T_1303_re <= _T_1302_re;
    _T_1303_im <= _T_1302_im;
    _T_1304_re <= _T_1303_re;
    _T_1304_im <= _T_1303_im;
    _T_1305_re <= _T_1304_re;
    _T_1305_im <= _T_1304_im;
    _T_1306_re <= _T_1305_re;
    _T_1306_im <= _T_1305_im;
    _T_1307_re <= _T_1306_re;
    _T_1307_im <= _T_1306_im;
    _T_1308_re <= _T_1307_re;
    _T_1308_im <= _T_1307_im;
    _T_1309_re <= _T_1308_re;
    _T_1309_im <= _T_1308_im;
    _T_1310_re <= _T_1309_re;
    _T_1310_im <= _T_1309_im;
    _T_1311_re <= _T_1310_re;
    _T_1311_im <= _T_1310_im;
    _T_1312_re <= _T_1311_re;
    _T_1312_im <= _T_1311_im;
    _T_1313_re <= _T_1312_re;
    _T_1313_im <= _T_1312_im;
    _T_1314_re <= _T_1313_re;
    _T_1314_im <= _T_1313_im;
    _T_1315_re <= _T_1314_re;
    _T_1315_im <= _T_1314_im;
    _T_1316_re <= _T_1315_re;
    _T_1316_im <= _T_1315_im;
    _T_1317_re <= _T_1316_re;
    _T_1317_im <= _T_1316_im;
    _T_1318_re <= _T_1317_re;
    _T_1318_im <= _T_1317_im;
    _T_1319_re <= _T_1318_re;
    _T_1319_im <= _T_1318_im;
    _T_1320_re <= _T_1319_re;
    _T_1320_im <= _T_1319_im;
    _T_1321_re <= _T_1320_re;
    _T_1321_im <= _T_1320_im;
    _T_1322_re <= _T_1321_re;
    _T_1322_im <= _T_1321_im;
    _T_1323_re <= _T_1322_re;
    _T_1323_im <= _T_1322_im;
    _T_1324_re <= _T_1323_re;
    _T_1324_im <= _T_1323_im;
    _T_1325_re <= _T_1324_re;
    _T_1325_im <= _T_1324_im;
    _T_1326_re <= _T_1325_re;
    _T_1326_im <= _T_1325_im;
    _T_1327_re <= _T_1326_re;
    _T_1327_im <= _T_1326_im;
    _T_1328_re <= _T_1327_re;
    _T_1328_im <= _T_1327_im;
    _T_1329_re <= _T_1328_re;
    _T_1329_im <= _T_1328_im;
    _T_1330_re <= _T_1329_re;
    _T_1330_im <= _T_1329_im;
    _T_1331_re <= _T_1330_re;
    _T_1331_im <= _T_1330_im;
    _T_1332_re <= _T_1331_re;
    _T_1332_im <= _T_1331_im;
    _T_1333_re <= _T_1332_re;
    _T_1333_im <= _T_1332_im;
    _T_1334_re <= _T_1333_re;
    _T_1334_im <= _T_1333_im;
    _T_1335_re <= _T_1334_re;
    _T_1335_im <= _T_1334_im;
    _T_1336_re <= _T_1335_re;
    _T_1336_im <= _T_1335_im;
    _T_1337_re <= _T_1336_re;
    _T_1337_im <= _T_1336_im;
    _T_1338_re <= _T_1337_re;
    _T_1338_im <= _T_1337_im;
    _T_1339_re <= _T_1338_re;
    _T_1339_im <= _T_1338_im;
    _T_1340_re <= _T_1339_re;
    _T_1340_im <= _T_1339_im;
    _T_1341_re <= _T_1340_re;
    _T_1341_im <= _T_1340_im;
    _T_1342_re <= _T_1341_re;
    _T_1342_im <= _T_1341_im;
    _T_1343_re <= _T_1342_re;
    _T_1343_im <= _T_1342_im;
    _T_1344_re <= _T_1343_re;
    _T_1344_im <= _T_1343_im;
    _T_1345_re <= _T_1344_re;
    _T_1345_im <= _T_1344_im;
    _T_1346_re <= _T_1345_re;
    _T_1346_im <= _T_1345_im;
    _T_1347_re <= _T_1346_re;
    _T_1347_im <= _T_1346_im;
    _T_1348_re <= _T_1347_re;
    _T_1348_im <= _T_1347_im;
    _T_1349_re <= _T_1348_re;
    _T_1349_im <= _T_1348_im;
    _T_1350_re <= _T_1349_re;
    _T_1350_im <= _T_1349_im;
    _T_1351_re <= _T_1350_re;
    _T_1351_im <= _T_1350_im;
    _T_1352_re <= _T_1351_re;
    _T_1352_im <= _T_1351_im;
    _T_1353_re <= _T_1352_re;
    _T_1353_im <= _T_1352_im;
    _T_1354_re <= _T_1353_re;
    _T_1354_im <= _T_1353_im;
    _T_1355_re <= _T_1354_re;
    _T_1355_im <= _T_1354_im;
    _T_1356_re <= _T_1355_re;
    _T_1356_im <= _T_1355_im;
    _T_1357_re <= _T_1356_re;
    _T_1357_im <= _T_1356_im;
    _T_1358_re <= _T_1357_re;
    _T_1358_im <= _T_1357_im;
    _T_1359_re <= _T_1358_re;
    _T_1359_im <= _T_1358_im;
    _T_1360_re <= _T_1359_re;
    _T_1360_im <= _T_1359_im;
    _T_1361_re <= _T_1360_re;
    _T_1361_im <= _T_1360_im;
    _T_1362_re <= _T_1361_re;
    _T_1362_im <= _T_1361_im;
    _T_1363_re <= _T_1362_re;
    _T_1363_im <= _T_1362_im;
    _T_1364_re <= _T_1363_re;
    _T_1364_im <= _T_1363_im;
    _T_1365_re <= _T_1364_re;
    _T_1365_im <= _T_1364_im;
    _T_1366_re <= _T_1365_re;
    _T_1366_im <= _T_1365_im;
    _T_1367_re <= _T_1366_re;
    _T_1367_im <= _T_1366_im;
    _T_1368_re <= _T_1367_re;
    _T_1368_im <= _T_1367_im;
    _T_1369_re <= _T_1368_re;
    _T_1369_im <= _T_1368_im;
    _T_1370_re <= _T_1369_re;
    _T_1370_im <= _T_1369_im;
    _T_1371_re <= _T_1370_re;
    _T_1371_im <= _T_1370_im;
    _T_1372_re <= _T_1371_re;
    _T_1372_im <= _T_1371_im;
    _T_1373_re <= _T_1372_re;
    _T_1373_im <= _T_1372_im;
    _T_1374_re <= _T_1373_re;
    _T_1374_im <= _T_1373_im;
    _T_1375_re <= _T_1374_re;
    _T_1375_im <= _T_1374_im;
    _T_1376_re <= _T_1375_re;
    _T_1376_im <= _T_1375_im;
    _T_1377_re <= _T_1376_re;
    _T_1377_im <= _T_1376_im;
    _T_1378_re <= _T_1377_re;
    _T_1378_im <= _T_1377_im;
    _T_1379_re <= _T_1378_re;
    _T_1379_im <= _T_1378_im;
    _T_1380_re <= _T_1379_re;
    _T_1380_im <= _T_1379_im;
    _T_1381_re <= _T_1380_re;
    _T_1381_im <= _T_1380_im;
    _T_1382_re <= _T_1381_re;
    _T_1382_im <= _T_1381_im;
    _T_1383_re <= _T_1382_re;
    _T_1383_im <= _T_1382_im;
    _T_1384_re <= _T_1383_re;
    _T_1384_im <= _T_1383_im;
    _T_1385_re <= _T_1384_re;
    _T_1385_im <= _T_1384_im;
    _T_1386_re <= _T_1385_re;
    _T_1386_im <= _T_1385_im;
    _T_1387_re <= _T_1386_re;
    _T_1387_im <= _T_1386_im;
    _T_1388_re <= _T_1387_re;
    _T_1388_im <= _T_1387_im;
    _T_1389_re <= _T_1388_re;
    _T_1389_im <= _T_1388_im;
    _T_1390_re <= _T_1389_re;
    _T_1390_im <= _T_1389_im;
    _T_1391_re <= _T_1390_re;
    _T_1391_im <= _T_1390_im;
    _T_1392_re <= _T_1391_re;
    _T_1392_im <= _T_1391_im;
    _T_1393_re <= _T_1392_re;
    _T_1393_im <= _T_1392_im;
    _T_1394_re <= _T_1393_re;
    _T_1394_im <= _T_1393_im;
    _T_1395_re <= _T_1394_re;
    _T_1395_im <= _T_1394_im;
    _T_1396_re <= _T_1395_re;
    _T_1396_im <= _T_1395_im;
    _T_1397_re <= _T_1396_re;
    _T_1397_im <= _T_1396_im;
    _T_1398_re <= _T_1397_re;
    _T_1398_im <= _T_1397_im;
    _T_1399_re <= _T_1398_re;
    _T_1399_im <= _T_1398_im;
    _T_1400_re <= _T_1399_re;
    _T_1400_im <= _T_1399_im;
    _T_1401_re <= _T_1400_re;
    _T_1401_im <= _T_1400_im;
    _T_1402_re <= _T_1401_re;
    _T_1402_im <= _T_1401_im;
    _T_1403_re <= _T_1402_re;
    _T_1403_im <= _T_1402_im;
    _T_1404_re <= _T_1403_re;
    _T_1404_im <= _T_1403_im;
    _T_1405_re <= _T_1404_re;
    _T_1405_im <= _T_1404_im;
    _T_1406_re <= _T_1405_re;
    _T_1406_im <= _T_1405_im;
    _T_1407_re <= _T_1406_re;
    _T_1407_im <= _T_1406_im;
    _T_1408_re <= _T_1407_re;
    _T_1408_im <= _T_1407_im;
    _T_1409_re <= _T_1408_re;
    _T_1409_im <= _T_1408_im;
    _T_1410_re <= _T_1409_re;
    _T_1410_im <= _T_1409_im;
    _T_1411_re <= _T_1410_re;
    _T_1411_im <= _T_1410_im;
    _T_1412_re <= _T_1411_re;
    _T_1412_im <= _T_1411_im;
    _T_1413_re <= _T_1412_re;
    _T_1413_im <= _T_1412_im;
    _T_1414_re <= _T_1413_re;
    _T_1414_im <= _T_1413_im;
    _T_1415_re <= _T_1414_re;
    _T_1415_im <= _T_1414_im;
    _T_1416_re <= _T_1415_re;
    _T_1416_im <= _T_1415_im;
    _T_1417_re <= _T_1416_re;
    _T_1417_im <= _T_1416_im;
    _T_1418_re <= _T_1417_re;
    _T_1418_im <= _T_1417_im;
    _T_1419_re <= _T_1418_re;
    _T_1419_im <= _T_1418_im;
    _T_1420_re <= _T_1419_re;
    _T_1420_im <= _T_1419_im;
    _T_1421_re <= _T_1420_re;
    _T_1421_im <= _T_1420_im;
    _T_1422_re <= _T_1421_re;
    _T_1422_im <= _T_1421_im;
    _T_1423_re <= _T_1422_re;
    _T_1423_im <= _T_1422_im;
    _T_1424_re <= _T_1423_re;
    _T_1424_im <= _T_1423_im;
    _T_1425_re <= _T_1424_re;
    _T_1425_im <= _T_1424_im;
    _T_1426_re <= _T_1425_re;
    _T_1426_im <= _T_1425_im;
    _T_1427_re <= _T_1426_re;
    _T_1427_im <= _T_1426_im;
    _T_1428_re <= _T_1427_re;
    _T_1428_im <= _T_1427_im;
    _T_1429_re <= _T_1428_re;
    _T_1429_im <= _T_1428_im;
    _T_1430_re <= _T_1429_re;
    _T_1430_im <= _T_1429_im;
    _T_1431_re <= _T_1430_re;
    _T_1431_im <= _T_1430_im;
    _T_1432_re <= _T_1431_re;
    _T_1432_im <= _T_1431_im;
    _T_1433_re <= _T_1432_re;
    _T_1433_im <= _T_1432_im;
    _T_1434_re <= _T_1433_re;
    _T_1434_im <= _T_1433_im;
    _T_1435_re <= _T_1434_re;
    _T_1435_im <= _T_1434_im;
    _T_1436_re <= _T_1435_re;
    _T_1436_im <= _T_1435_im;
    _T_1437_re <= _T_1436_re;
    _T_1437_im <= _T_1436_im;
    _T_1438_re <= _T_1437_re;
    _T_1438_im <= _T_1437_im;
    _T_1439_re <= _T_1438_re;
    _T_1439_im <= _T_1438_im;
    _T_1440_re <= _T_1439_re;
    _T_1440_im <= _T_1439_im;
    _T_1441_re <= _T_1440_re;
    _T_1441_im <= _T_1440_im;
    _T_1442_re <= _T_1441_re;
    _T_1442_im <= _T_1441_im;
    _T_1443_re <= _T_1442_re;
    _T_1443_im <= _T_1442_im;
    _T_1444_re <= _T_1443_re;
    _T_1444_im <= _T_1443_im;
    _T_1445_re <= _T_1444_re;
    _T_1445_im <= _T_1444_im;
    _T_1446_re <= _T_1445_re;
    _T_1446_im <= _T_1445_im;
    _T_1447_re <= _T_1446_re;
    _T_1447_im <= _T_1446_im;
    _T_1448_re <= _T_1447_re;
    _T_1448_im <= _T_1447_im;
    _T_1449_re <= _T_1448_re;
    _T_1449_im <= _T_1448_im;
    _T_1450_re <= _T_1449_re;
    _T_1450_im <= _T_1449_im;
    _T_1451_re <= _T_1450_re;
    _T_1451_im <= _T_1450_im;
    _T_1452_re <= _T_1451_re;
    _T_1452_im <= _T_1451_im;
    _T_1453_re <= _T_1452_re;
    _T_1453_im <= _T_1452_im;
    _T_1454_re <= _T_1453_re;
    _T_1454_im <= _T_1453_im;
    _T_1455_re <= _T_1454_re;
    _T_1455_im <= _T_1454_im;
    _T_1456_re <= _T_1455_re;
    _T_1456_im <= _T_1455_im;
    _T_1457_re <= _T_1456_re;
    _T_1457_im <= _T_1456_im;
    _T_1458_re <= _T_1457_re;
    _T_1458_im <= _T_1457_im;
    _T_1459_re <= _T_1458_re;
    _T_1459_im <= _T_1458_im;
    _T_1460_re <= _T_1459_re;
    _T_1460_im <= _T_1459_im;
    _T_1461_re <= _T_1460_re;
    _T_1461_im <= _T_1460_im;
    _T_1462_re <= _T_1461_re;
    _T_1462_im <= _T_1461_im;
    _T_1463_re <= _T_1462_re;
    _T_1463_im <= _T_1462_im;
    _T_1464_re <= _T_1463_re;
    _T_1464_im <= _T_1463_im;
    _T_1465_re <= _T_1464_re;
    _T_1465_im <= _T_1464_im;
    _T_1466_re <= _T_1465_re;
    _T_1466_im <= _T_1465_im;
    _T_1467_re <= _T_1466_re;
    _T_1467_im <= _T_1466_im;
    _T_1468_re <= _T_1467_re;
    _T_1468_im <= _T_1467_im;
    _T_1469_re <= _T_1468_re;
    _T_1469_im <= _T_1468_im;
    _T_1470_re <= _T_1469_re;
    _T_1470_im <= _T_1469_im;
    _T_1471_re <= _T_1470_re;
    _T_1471_im <= _T_1470_im;
    _T_1472_re <= _T_1471_re;
    _T_1472_im <= _T_1471_im;
    _T_1473_re <= _T_1472_re;
    _T_1473_im <= _T_1472_im;
    _T_1474_re <= _T_1473_re;
    _T_1474_im <= _T_1473_im;
    _T_1475_re <= _T_1474_re;
    _T_1475_im <= _T_1474_im;
    _T_1476_re <= _T_1475_re;
    _T_1476_im <= _T_1475_im;
    _T_1477_re <= _T_1476_re;
    _T_1477_im <= _T_1476_im;
    _T_1478_re <= _T_1477_re;
    _T_1478_im <= _T_1477_im;
    _T_1479_re <= _T_1478_re;
    _T_1479_im <= _T_1478_im;
    _T_1480_re <= _T_1479_re;
    _T_1480_im <= _T_1479_im;
    _T_1481_re <= _T_1480_re;
    _T_1481_im <= _T_1480_im;
    _T_1482_re <= _T_1481_re;
    _T_1482_im <= _T_1481_im;
    _T_1483_re <= _T_1482_re;
    _T_1483_im <= _T_1482_im;
    _T_1484_re <= _T_1483_re;
    _T_1484_im <= _T_1483_im;
    _T_1485_re <= _T_1484_re;
    _T_1485_im <= _T_1484_im;
    _T_1486_re <= _T_1485_re;
    _T_1486_im <= _T_1485_im;
    _T_1487_re <= _T_1486_re;
    _T_1487_im <= _T_1486_im;
    _T_1488_re <= _T_1487_re;
    _T_1488_im <= _T_1487_im;
    _T_1489_re <= _T_1488_re;
    _T_1489_im <= _T_1488_im;
    _T_1490_re <= _T_1489_re;
    _T_1490_im <= _T_1489_im;
    _T_1491_re <= _T_1490_re;
    _T_1491_im <= _T_1490_im;
    _T_1492_re <= _T_1491_re;
    _T_1492_im <= _T_1491_im;
    _T_1493_re <= _T_1492_re;
    _T_1493_im <= _T_1492_im;
    _T_1494_re <= _T_1493_re;
    _T_1494_im <= _T_1493_im;
    _T_1495_re <= _T_1494_re;
    _T_1495_im <= _T_1494_im;
    _T_1496_re <= _T_1495_re;
    _T_1496_im <= _T_1495_im;
    _T_1497_re <= _T_1496_re;
    _T_1497_im <= _T_1496_im;
    _T_1498_re <= _T_1497_re;
    _T_1498_im <= _T_1497_im;
    _T_1499_re <= _T_1498_re;
    _T_1499_im <= _T_1498_im;
    _T_1500_re <= _T_1499_re;
    _T_1500_im <= _T_1499_im;
    _T_1501_re <= _T_1500_re;
    _T_1501_im <= _T_1500_im;
    _T_1502_re <= _T_1501_re;
    _T_1502_im <= _T_1501_im;
    _T_1503_re <= _T_1502_re;
    _T_1503_im <= _T_1502_im;
    _T_1504_re <= _T_1503_re;
    _T_1504_im <= _T_1503_im;
    _T_1505_re <= _T_1504_re;
    _T_1505_im <= _T_1504_im;
    _T_1506_re <= _T_1505_re;
    _T_1506_im <= _T_1505_im;
    _T_1507_re <= _T_1506_re;
    _T_1507_im <= _T_1506_im;
    _T_1508_re <= _T_1507_re;
    _T_1508_im <= _T_1507_im;
    _T_1509_re <= _T_1508_re;
    _T_1509_im <= _T_1508_im;
    _T_1510_re <= _T_1509_re;
    _T_1510_im <= _T_1509_im;
    _T_1511_re <= _T_1510_re;
    _T_1511_im <= _T_1510_im;
    _T_1512_re <= _T_1511_re;
    _T_1512_im <= _T_1511_im;
    _T_1513_re <= _T_1512_re;
    _T_1513_im <= _T_1512_im;
    _T_1514_re <= _T_1513_re;
    _T_1514_im <= _T_1513_im;
    _T_1515_re <= _T_1514_re;
    _T_1515_im <= _T_1514_im;
    _T_1516_re <= _T_1515_re;
    _T_1516_im <= _T_1515_im;
    _T_1517_re <= _T_1516_re;
    _T_1517_im <= _T_1516_im;
    _T_1518_re <= _T_1517_re;
    _T_1518_im <= _T_1517_im;
    _T_1519_re <= _T_1518_re;
    _T_1519_im <= _T_1518_im;
    _T_1520_re <= _T_1519_re;
    _T_1520_im <= _T_1519_im;
    _T_1521_re <= _T_1520_re;
    _T_1521_im <= _T_1520_im;
    _T_1522_re <= _T_1521_re;
    _T_1522_im <= _T_1521_im;
    _T_1523_re <= _T_1522_re;
    _T_1523_im <= _T_1522_im;
    _T_1524_re <= _T_1523_re;
    _T_1524_im <= _T_1523_im;
    _T_1525_re <= _T_1524_re;
    _T_1525_im <= _T_1524_im;
    _T_1526_re <= _T_1525_re;
    _T_1526_im <= _T_1525_im;
    _T_1527_re <= _T_1526_re;
    _T_1527_im <= _T_1526_im;
    _T_1528_re <= _T_1527_re;
    _T_1528_im <= _T_1527_im;
    _T_1529_re <= _T_1528_re;
    _T_1529_im <= _T_1528_im;
    _T_1530_re <= _T_1529_re;
    _T_1530_im <= _T_1529_im;
    _T_1531_re <= _T_1530_re;
    _T_1531_im <= _T_1530_im;
    _T_1532_re <= _T_1531_re;
    _T_1532_im <= _T_1531_im;
    _T_1533_re <= _T_1532_re;
    _T_1533_im <= _T_1532_im;
    _T_1534_re <= _T_1533_re;
    _T_1534_im <= _T_1533_im;
    _T_1535_re <= _T_1534_re;
    _T_1535_im <= _T_1534_im;
    _T_1536_re <= _T_1535_re;
    _T_1536_im <= _T_1535_im;
    _T_1537_re <= _T_1536_re;
    _T_1537_im <= _T_1536_im;
    _T_1538_re <= _T_1537_re;
    _T_1538_im <= _T_1537_im;
    _T_1539_re <= _T_1538_re;
    _T_1539_im <= _T_1538_im;
    _T_1540_re <= _T_1539_re;
    _T_1540_im <= _T_1539_im;
    _T_1541_re <= _T_1540_re;
    _T_1541_im <= _T_1540_im;
    _T_1542_re <= _T_1541_re;
    _T_1542_im <= _T_1541_im;
    _T_1543_re <= _T_1542_re;
    _T_1543_im <= _T_1542_im;
    _T_1544_re <= _T_1543_re;
    _T_1544_im <= _T_1543_im;
    _T_1545_re <= _T_1544_re;
    _T_1545_im <= _T_1544_im;
    _T_1546_re <= _T_1545_re;
    _T_1546_im <= _T_1545_im;
    _T_1547_re <= _T_1546_re;
    _T_1547_im <= _T_1546_im;
    _T_1548_re <= _T_1547_re;
    _T_1548_im <= _T_1547_im;
    _T_1549_re <= _T_1548_re;
    _T_1549_im <= _T_1548_im;
    _T_1550_re <= _T_1549_re;
    _T_1550_im <= _T_1549_im;
    _T_1551_re <= _T_1550_re;
    _T_1551_im <= _T_1550_im;
    _T_1552_re <= _T_1551_re;
    _T_1552_im <= _T_1551_im;
    _T_1553_re <= _T_1552_re;
    _T_1553_im <= _T_1552_im;
    _T_1554_re <= _T_1553_re;
    _T_1554_im <= _T_1553_im;
    _T_1555_re <= _T_1554_re;
    _T_1555_im <= _T_1554_im;
    _T_1556_re <= _T_1555_re;
    _T_1556_im <= _T_1555_im;
    _T_1557_re <= _T_1556_re;
    _T_1557_im <= _T_1556_im;
    _T_1558_re <= _T_1557_re;
    _T_1558_im <= _T_1557_im;
    _T_1559_re <= _T_1558_re;
    _T_1559_im <= _T_1558_im;
    _T_1560_re <= _T_1559_re;
    _T_1560_im <= _T_1559_im;
    _T_1561_re <= _T_1560_re;
    _T_1561_im <= _T_1560_im;
    _T_1562_re <= _T_1561_re;
    _T_1562_im <= _T_1561_im;
    _T_1563_re <= _T_1562_re;
    _T_1563_im <= _T_1562_im;
    _T_1564_re <= _T_1563_re;
    _T_1564_im <= _T_1563_im;
    _T_1565_re <= _T_1564_re;
    _T_1565_im <= _T_1564_im;
    _T_1566_re <= _T_1565_re;
    _T_1566_im <= _T_1565_im;
    _T_1567_re <= _T_1566_re;
    _T_1567_im <= _T_1566_im;
    _T_1568_re <= _T_1567_re;
    _T_1568_im <= _T_1567_im;
    _T_1569_re <= _T_1568_re;
    _T_1569_im <= _T_1568_im;
    _T_1570_re <= _T_1569_re;
    _T_1570_im <= _T_1569_im;
    _T_1571_re <= _T_1570_re;
    _T_1571_im <= _T_1570_im;
    _T_1572_re <= _T_1571_re;
    _T_1572_im <= _T_1571_im;
    _T_1573_re <= _T_1572_re;
    _T_1573_im <= _T_1572_im;
    _T_1574_re <= _T_1573_re;
    _T_1574_im <= _T_1573_im;
    _T_1575_re <= _T_1574_re;
    _T_1575_im <= _T_1574_im;
    _T_1576_re <= _T_1575_re;
    _T_1576_im <= _T_1575_im;
    _T_1577_re <= _T_1576_re;
    _T_1577_im <= _T_1576_im;
    _T_1578_re <= _T_1577_re;
    _T_1578_im <= _T_1577_im;
    _T_1579_re <= _T_1578_re;
    _T_1579_im <= _T_1578_im;
    _T_1580_re <= _T_1579_re;
    _T_1580_im <= _T_1579_im;
    _T_1581_re <= _T_1580_re;
    _T_1581_im <= _T_1580_im;
    _T_1582_re <= _T_1581_re;
    _T_1582_im <= _T_1581_im;
    _T_1583_re <= _T_1582_re;
    _T_1583_im <= _T_1582_im;
    _T_1584_re <= _T_1583_re;
    _T_1584_im <= _T_1583_im;
    _T_1585_re <= _T_1584_re;
    _T_1585_im <= _T_1584_im;
    _T_1586_re <= _T_1585_re;
    _T_1586_im <= _T_1585_im;
    _T_1587_re <= _T_1586_re;
    _T_1587_im <= _T_1586_im;
    _T_1588_re <= _T_1587_re;
    _T_1588_im <= _T_1587_im;
    _T_1589_re <= _T_1588_re;
    _T_1589_im <= _T_1588_im;
    _T_1590_re <= _T_1589_re;
    _T_1590_im <= _T_1589_im;
    _T_1591_re <= _T_1590_re;
    _T_1591_im <= _T_1590_im;
    _T_1592_re <= _T_1591_re;
    _T_1592_im <= _T_1591_im;
    _T_1593_re <= _T_1592_re;
    _T_1593_im <= _T_1592_im;
    _T_1594_re <= _T_1593_re;
    _T_1594_im <= _T_1593_im;
    _T_1595_re <= _T_1594_re;
    _T_1595_im <= _T_1594_im;
    _T_1596_re <= _T_1595_re;
    _T_1596_im <= _T_1595_im;
    _T_1597_re <= _T_1596_re;
    _T_1597_im <= _T_1596_im;
    _T_1598_re <= _T_1597_re;
    _T_1598_im <= _T_1597_im;
    _T_1599_re <= _T_1598_re;
    _T_1599_im <= _T_1598_im;
    _T_1600_re <= _T_1599_re;
    _T_1600_im <= _T_1599_im;
    _T_1601_re <= _T_1600_re;
    _T_1601_im <= _T_1600_im;
    _T_1602_re <= _T_1601_re;
    _T_1602_im <= _T_1601_im;
    _T_1603_re <= _T_1602_re;
    _T_1603_im <= _T_1602_im;
    _T_1604_re <= _T_1603_re;
    _T_1604_im <= _T_1603_im;
    _T_1605_re <= _T_1604_re;
    _T_1605_im <= _T_1604_im;
    _T_1606_re <= _T_1605_re;
    _T_1606_im <= _T_1605_im;
    _T_1607_re <= _T_1606_re;
    _T_1607_im <= _T_1606_im;
    _T_1608_re <= _T_1607_re;
    _T_1608_im <= _T_1607_im;
    _T_1609_re <= _T_1608_re;
    _T_1609_im <= _T_1608_im;
    _T_1610_re <= _T_1609_re;
    _T_1610_im <= _T_1609_im;
    _T_1611_re <= _T_1610_re;
    _T_1611_im <= _T_1610_im;
    _T_1612_re <= _T_1611_re;
    _T_1612_im <= _T_1611_im;
    _T_1613_re <= _T_1612_re;
    _T_1613_im <= _T_1612_im;
    _T_1614_re <= _T_1613_re;
    _T_1614_im <= _T_1613_im;
    _T_1615_re <= _T_1614_re;
    _T_1615_im <= _T_1614_im;
    _T_1616_re <= _T_1615_re;
    _T_1616_im <= _T_1615_im;
    _T_1617_re <= _T_1616_re;
    _T_1617_im <= _T_1616_im;
    _T_1618_re <= _T_1617_re;
    _T_1618_im <= _T_1617_im;
    _T_1619_re <= _T_1618_re;
    _T_1619_im <= _T_1618_im;
    _T_1620_re <= _T_1619_re;
    _T_1620_im <= _T_1619_im;
    _T_1621_re <= _T_1620_re;
    _T_1621_im <= _T_1620_im;
    _T_1622_re <= _T_1621_re;
    _T_1622_im <= _T_1621_im;
    _T_1623_re <= _T_1622_re;
    _T_1623_im <= _T_1622_im;
    _T_1624_re <= _T_1623_re;
    _T_1624_im <= _T_1623_im;
    _T_1625_re <= _T_1624_re;
    _T_1625_im <= _T_1624_im;
    _T_1626_re <= _T_1625_re;
    _T_1626_im <= _T_1625_im;
    _T_1627_re <= _T_1626_re;
    _T_1627_im <= _T_1626_im;
    _T_1628_re <= _T_1627_re;
    _T_1628_im <= _T_1627_im;
    _T_1629_re <= _T_1628_re;
    _T_1629_im <= _T_1628_im;
    _T_1630_re <= _T_1629_re;
    _T_1630_im <= _T_1629_im;
    _T_1631_re <= _T_1630_re;
    _T_1631_im <= _T_1630_im;
    _T_1632_re <= _T_1631_re;
    _T_1632_im <= _T_1631_im;
    _T_1633_re <= _T_1632_re;
    _T_1633_im <= _T_1632_im;
    _T_1634_re <= _T_1633_re;
    _T_1634_im <= _T_1633_im;
    _T_1635_re <= _T_1634_re;
    _T_1635_im <= _T_1634_im;
    _T_1636_re <= _T_1635_re;
    _T_1636_im <= _T_1635_im;
    _T_1637_re <= _T_1636_re;
    _T_1637_im <= _T_1636_im;
    _T_1638_re <= _T_1637_re;
    _T_1638_im <= _T_1637_im;
    _T_1639_re <= _T_1638_re;
    _T_1639_im <= _T_1638_im;
    _T_1640_re <= _T_1639_re;
    _T_1640_im <= _T_1639_im;
    _T_1641_re <= _T_1640_re;
    _T_1641_im <= _T_1640_im;
    _T_1642_re <= _T_1641_re;
    _T_1642_im <= _T_1641_im;
    _T_1643_re <= _T_1642_re;
    _T_1643_im <= _T_1642_im;
    _T_1644_re <= _T_1643_re;
    _T_1644_im <= _T_1643_im;
    _T_1645_re <= _T_1644_re;
    _T_1645_im <= _T_1644_im;
    _T_1646_re <= _T_1645_re;
    _T_1646_im <= _T_1645_im;
    _T_1647_re <= _T_1646_re;
    _T_1647_im <= _T_1646_im;
    _T_1648_re <= _T_1647_re;
    _T_1648_im <= _T_1647_im;
    _T_1649_re <= _T_1648_re;
    _T_1649_im <= _T_1648_im;
    _T_1650_re <= _T_1649_re;
    _T_1650_im <= _T_1649_im;
    _T_1651_re <= _T_1650_re;
    _T_1651_im <= _T_1650_im;
    _T_1652_re <= _T_1651_re;
    _T_1652_im <= _T_1651_im;
    _T_1653_re <= _T_1652_re;
    _T_1653_im <= _T_1652_im;
    _T_1654_re <= _T_1653_re;
    _T_1654_im <= _T_1653_im;
    _T_1655_re <= _T_1654_re;
    _T_1655_im <= _T_1654_im;
    _T_1656_re <= _T_1655_re;
    _T_1656_im <= _T_1655_im;
    _T_1657_re <= _T_1656_re;
    _T_1657_im <= _T_1656_im;
    _T_1658_re <= _T_1657_re;
    _T_1658_im <= _T_1657_im;
    _T_1659_re <= _T_1658_re;
    _T_1659_im <= _T_1658_im;
    _T_1660_re <= _T_1659_re;
    _T_1660_im <= _T_1659_im;
    _T_1661_re <= _T_1660_re;
    _T_1661_im <= _T_1660_im;
    _T_1662_re <= _T_1661_re;
    _T_1662_im <= _T_1661_im;
    _T_1663_re <= _T_1662_re;
    _T_1663_im <= _T_1662_im;
    _T_1664_re <= _T_1663_re;
    _T_1664_im <= _T_1663_im;
    _T_1665_re <= _T_1664_re;
    _T_1665_im <= _T_1664_im;
    _T_1666_re <= _T_1665_re;
    _T_1666_im <= _T_1665_im;
    _T_1667_re <= _T_1666_re;
    _T_1667_im <= _T_1666_im;
    _T_1668_re <= _T_1667_re;
    _T_1668_im <= _T_1667_im;
    _T_1669_re <= _T_1668_re;
    _T_1669_im <= _T_1668_im;
    _T_1670_re <= _T_1669_re;
    _T_1670_im <= _T_1669_im;
    _T_1671_re <= _T_1670_re;
    _T_1671_im <= _T_1670_im;
    _T_1672_re <= _T_1671_re;
    _T_1672_im <= _T_1671_im;
    _T_1673_re <= _T_1672_re;
    _T_1673_im <= _T_1672_im;
    _T_1674_re <= _T_1673_re;
    _T_1674_im <= _T_1673_im;
    _T_1675_re <= _T_1674_re;
    _T_1675_im <= _T_1674_im;
    _T_1676_re <= _T_1675_re;
    _T_1676_im <= _T_1675_im;
    _T_1677_re <= _T_1676_re;
    _T_1677_im <= _T_1676_im;
    _T_1678_re <= _T_1677_re;
    _T_1678_im <= _T_1677_im;
    _T_1679_re <= _T_1678_re;
    _T_1679_im <= _T_1678_im;
    _T_1680_re <= _T_1679_re;
    _T_1680_im <= _T_1679_im;
    _T_1681_re <= _T_1680_re;
    _T_1681_im <= _T_1680_im;
    _T_1682_re <= _T_1681_re;
    _T_1682_im <= _T_1681_im;
    _T_1683_re <= _T_1682_re;
    _T_1683_im <= _T_1682_im;
    _T_1684_re <= _T_1683_re;
    _T_1684_im <= _T_1683_im;
    _T_1685_re <= _T_1684_re;
    _T_1685_im <= _T_1684_im;
    _T_1686_re <= _T_1685_re;
    _T_1686_im <= _T_1685_im;
    _T_1687_re <= _T_1686_re;
    _T_1687_im <= _T_1686_im;
    _T_1688_re <= _T_1687_re;
    _T_1688_im <= _T_1687_im;
    _T_1689_re <= _T_1688_re;
    _T_1689_im <= _T_1688_im;
    _T_1690_re <= _T_1689_re;
    _T_1690_im <= _T_1689_im;
    _T_1691_re <= _T_1690_re;
    _T_1691_im <= _T_1690_im;
    _T_1692_re <= _T_1691_re;
    _T_1692_im <= _T_1691_im;
    _T_1693_re <= _T_1692_re;
    _T_1693_im <= _T_1692_im;
    _T_1694_re <= _T_1693_re;
    _T_1694_im <= _T_1693_im;
    _T_1695_re <= _T_1694_re;
    _T_1695_im <= _T_1694_im;
    _T_1696_re <= _T_1695_re;
    _T_1696_im <= _T_1695_im;
    _T_1697_re <= _T_1696_re;
    _T_1697_im <= _T_1696_im;
    _T_1698_re <= _T_1697_re;
    _T_1698_im <= _T_1697_im;
    _T_1699_re <= _T_1698_re;
    _T_1699_im <= _T_1698_im;
    _T_1700_re <= _T_1699_re;
    _T_1700_im <= _T_1699_im;
    _T_1701_re <= _T_1700_re;
    _T_1701_im <= _T_1700_im;
    _T_1702_re <= _T_1701_re;
    _T_1702_im <= _T_1701_im;
    _T_1703_re <= _T_1702_re;
    _T_1703_im <= _T_1702_im;
    _T_1704_re <= _T_1703_re;
    _T_1704_im <= _T_1703_im;
    _T_1705_re <= _T_1704_re;
    _T_1705_im <= _T_1704_im;
    _T_1706_re <= _T_1705_re;
    _T_1706_im <= _T_1705_im;
    _T_1707_re <= _T_1706_re;
    _T_1707_im <= _T_1706_im;
    _T_1708_re <= _T_1707_re;
    _T_1708_im <= _T_1707_im;
    _T_1709_re <= _T_1708_re;
    _T_1709_im <= _T_1708_im;
    _T_1710_re <= _T_1709_re;
    _T_1710_im <= _T_1709_im;
    _T_1711_re <= _T_1710_re;
    _T_1711_im <= _T_1710_im;
    _T_1712_re <= _T_1711_re;
    _T_1712_im <= _T_1711_im;
    _T_1713_re <= _T_1712_re;
    _T_1713_im <= _T_1712_im;
    _T_1714_re <= _T_1713_re;
    _T_1714_im <= _T_1713_im;
    _T_1715_re <= _T_1714_re;
    _T_1715_im <= _T_1714_im;
    _T_1716_re <= _T_1715_re;
    _T_1716_im <= _T_1715_im;
    _T_1717_re <= _T_1716_re;
    _T_1717_im <= _T_1716_im;
    _T_1718_re <= _T_1717_re;
    _T_1718_im <= _T_1717_im;
    _T_1728_re <= Switch_io_out1_re;
    _T_1728_im <= Switch_io_out1_im;
    _T_1729_re <= _T_1728_re;
    _T_1729_im <= _T_1728_im;
    _T_1730_re <= _T_1729_re;
    _T_1730_im <= _T_1729_im;
    _T_1731_re <= _T_1730_re;
    _T_1731_im <= _T_1730_im;
    _T_1732_re <= _T_1731_re;
    _T_1732_im <= _T_1731_im;
    _T_1733_re <= _T_1732_re;
    _T_1733_im <= _T_1732_im;
    _T_1734_re <= _T_1733_re;
    _T_1734_im <= _T_1733_im;
    _T_1735_re <= _T_1734_re;
    _T_1735_im <= _T_1734_im;
    _T_1736_re <= _T_1735_re;
    _T_1736_im <= _T_1735_im;
    _T_1737_re <= _T_1736_re;
    _T_1737_im <= _T_1736_im;
    _T_1738_re <= _T_1737_re;
    _T_1738_im <= _T_1737_im;
    _T_1739_re <= _T_1738_re;
    _T_1739_im <= _T_1738_im;
    _T_1740_re <= _T_1739_re;
    _T_1740_im <= _T_1739_im;
    _T_1741_re <= _T_1740_re;
    _T_1741_im <= _T_1740_im;
    _T_1742_re <= _T_1741_re;
    _T_1742_im <= _T_1741_im;
    _T_1743_re <= _T_1742_re;
    _T_1743_im <= _T_1742_im;
    _T_1744_re <= _T_1743_re;
    _T_1744_im <= _T_1743_im;
    _T_1745_re <= _T_1744_re;
    _T_1745_im <= _T_1744_im;
    _T_1746_re <= _T_1745_re;
    _T_1746_im <= _T_1745_im;
    _T_1747_re <= _T_1746_re;
    _T_1747_im <= _T_1746_im;
    _T_1748_re <= _T_1747_re;
    _T_1748_im <= _T_1747_im;
    _T_1749_re <= _T_1748_re;
    _T_1749_im <= _T_1748_im;
    _T_1750_re <= _T_1749_re;
    _T_1750_im <= _T_1749_im;
    _T_1751_re <= _T_1750_re;
    _T_1751_im <= _T_1750_im;
    _T_1752_re <= _T_1751_re;
    _T_1752_im <= _T_1751_im;
    _T_1753_re <= _T_1752_re;
    _T_1753_im <= _T_1752_im;
    _T_1754_re <= _T_1753_re;
    _T_1754_im <= _T_1753_im;
    _T_1755_re <= _T_1754_re;
    _T_1755_im <= _T_1754_im;
    _T_1756_re <= _T_1755_re;
    _T_1756_im <= _T_1755_im;
    _T_1757_re <= _T_1756_re;
    _T_1757_im <= _T_1756_im;
    _T_1758_re <= _T_1757_re;
    _T_1758_im <= _T_1757_im;
    _T_1759_re <= _T_1758_re;
    _T_1759_im <= _T_1758_im;
    _T_1760_re <= _T_1759_re;
    _T_1760_im <= _T_1759_im;
    _T_1761_re <= _T_1760_re;
    _T_1761_im <= _T_1760_im;
    _T_1762_re <= _T_1761_re;
    _T_1762_im <= _T_1761_im;
    _T_1763_re <= _T_1762_re;
    _T_1763_im <= _T_1762_im;
    _T_1764_re <= _T_1763_re;
    _T_1764_im <= _T_1763_im;
    _T_1765_re <= _T_1764_re;
    _T_1765_im <= _T_1764_im;
    _T_1766_re <= _T_1765_re;
    _T_1766_im <= _T_1765_im;
    _T_1767_re <= _T_1766_re;
    _T_1767_im <= _T_1766_im;
    _T_1768_re <= _T_1767_re;
    _T_1768_im <= _T_1767_im;
    _T_1769_re <= _T_1768_re;
    _T_1769_im <= _T_1768_im;
    _T_1770_re <= _T_1769_re;
    _T_1770_im <= _T_1769_im;
    _T_1771_re <= _T_1770_re;
    _T_1771_im <= _T_1770_im;
    _T_1772_re <= _T_1771_re;
    _T_1772_im <= _T_1771_im;
    _T_1773_re <= _T_1772_re;
    _T_1773_im <= _T_1772_im;
    _T_1774_re <= _T_1773_re;
    _T_1774_im <= _T_1773_im;
    _T_1775_re <= _T_1774_re;
    _T_1775_im <= _T_1774_im;
    _T_1776_re <= _T_1775_re;
    _T_1776_im <= _T_1775_im;
    _T_1777_re <= _T_1776_re;
    _T_1777_im <= _T_1776_im;
    _T_1778_re <= _T_1777_re;
    _T_1778_im <= _T_1777_im;
    _T_1779_re <= _T_1778_re;
    _T_1779_im <= _T_1778_im;
    _T_1780_re <= _T_1779_re;
    _T_1780_im <= _T_1779_im;
    _T_1781_re <= _T_1780_re;
    _T_1781_im <= _T_1780_im;
    _T_1782_re <= _T_1781_re;
    _T_1782_im <= _T_1781_im;
    _T_1783_re <= _T_1782_re;
    _T_1783_im <= _T_1782_im;
    _T_1784_re <= _T_1783_re;
    _T_1784_im <= _T_1783_im;
    _T_1785_re <= _T_1784_re;
    _T_1785_im <= _T_1784_im;
    _T_1786_re <= _T_1785_re;
    _T_1786_im <= _T_1785_im;
    _T_1787_re <= _T_1786_re;
    _T_1787_im <= _T_1786_im;
    _T_1788_re <= _T_1787_re;
    _T_1788_im <= _T_1787_im;
    _T_1789_re <= _T_1788_re;
    _T_1789_im <= _T_1788_im;
    _T_1790_re <= _T_1789_re;
    _T_1790_im <= _T_1789_im;
    _T_1791_re <= _T_1790_re;
    _T_1791_im <= _T_1790_im;
    _T_1792_re <= _T_1791_re;
    _T_1792_im <= _T_1791_im;
    _T_1793_re <= _T_1792_re;
    _T_1793_im <= _T_1792_im;
    _T_1794_re <= _T_1793_re;
    _T_1794_im <= _T_1793_im;
    _T_1795_re <= _T_1794_re;
    _T_1795_im <= _T_1794_im;
    _T_1796_re <= _T_1795_re;
    _T_1796_im <= _T_1795_im;
    _T_1797_re <= _T_1796_re;
    _T_1797_im <= _T_1796_im;
    _T_1798_re <= _T_1797_re;
    _T_1798_im <= _T_1797_im;
    _T_1799_re <= _T_1798_re;
    _T_1799_im <= _T_1798_im;
    _T_1800_re <= _T_1799_re;
    _T_1800_im <= _T_1799_im;
    _T_1801_re <= _T_1800_re;
    _T_1801_im <= _T_1800_im;
    _T_1802_re <= _T_1801_re;
    _T_1802_im <= _T_1801_im;
    _T_1803_re <= _T_1802_re;
    _T_1803_im <= _T_1802_im;
    _T_1804_re <= _T_1803_re;
    _T_1804_im <= _T_1803_im;
    _T_1805_re <= _T_1804_re;
    _T_1805_im <= _T_1804_im;
    _T_1806_re <= _T_1805_re;
    _T_1806_im <= _T_1805_im;
    _T_1807_re <= _T_1806_re;
    _T_1807_im <= _T_1806_im;
    _T_1808_re <= _T_1807_re;
    _T_1808_im <= _T_1807_im;
    _T_1809_re <= _T_1808_re;
    _T_1809_im <= _T_1808_im;
    _T_1810_re <= _T_1809_re;
    _T_1810_im <= _T_1809_im;
    _T_1811_re <= _T_1810_re;
    _T_1811_im <= _T_1810_im;
    _T_1812_re <= _T_1811_re;
    _T_1812_im <= _T_1811_im;
    _T_1813_re <= _T_1812_re;
    _T_1813_im <= _T_1812_im;
    _T_1814_re <= _T_1813_re;
    _T_1814_im <= _T_1813_im;
    _T_1815_re <= _T_1814_re;
    _T_1815_im <= _T_1814_im;
    _T_1816_re <= _T_1815_re;
    _T_1816_im <= _T_1815_im;
    _T_1817_re <= _T_1816_re;
    _T_1817_im <= _T_1816_im;
    _T_1818_re <= _T_1817_re;
    _T_1818_im <= _T_1817_im;
    _T_1819_re <= _T_1818_re;
    _T_1819_im <= _T_1818_im;
    _T_1820_re <= _T_1819_re;
    _T_1820_im <= _T_1819_im;
    _T_1821_re <= _T_1820_re;
    _T_1821_im <= _T_1820_im;
    _T_1822_re <= _T_1821_re;
    _T_1822_im <= _T_1821_im;
    _T_1823_re <= _T_1822_re;
    _T_1823_im <= _T_1822_im;
    _T_1824_re <= _T_1823_re;
    _T_1824_im <= _T_1823_im;
    _T_1825_re <= _T_1824_re;
    _T_1825_im <= _T_1824_im;
    _T_1826_re <= _T_1825_re;
    _T_1826_im <= _T_1825_im;
    _T_1827_re <= _T_1826_re;
    _T_1827_im <= _T_1826_im;
    _T_1828_re <= _T_1827_re;
    _T_1828_im <= _T_1827_im;
    _T_1829_re <= _T_1828_re;
    _T_1829_im <= _T_1828_im;
    _T_1830_re <= _T_1829_re;
    _T_1830_im <= _T_1829_im;
    _T_1831_re <= _T_1830_re;
    _T_1831_im <= _T_1830_im;
    _T_1832_re <= _T_1831_re;
    _T_1832_im <= _T_1831_im;
    _T_1833_re <= _T_1832_re;
    _T_1833_im <= _T_1832_im;
    _T_1834_re <= _T_1833_re;
    _T_1834_im <= _T_1833_im;
    _T_1835_re <= _T_1834_re;
    _T_1835_im <= _T_1834_im;
    _T_1836_re <= _T_1835_re;
    _T_1836_im <= _T_1835_im;
    _T_1837_re <= _T_1836_re;
    _T_1837_im <= _T_1836_im;
    _T_1838_re <= _T_1837_re;
    _T_1838_im <= _T_1837_im;
    _T_1839_re <= _T_1838_re;
    _T_1839_im <= _T_1838_im;
    _T_1840_re <= _T_1839_re;
    _T_1840_im <= _T_1839_im;
    _T_1841_re <= _T_1840_re;
    _T_1841_im <= _T_1840_im;
    _T_1842_re <= _T_1841_re;
    _T_1842_im <= _T_1841_im;
    _T_1843_re <= _T_1842_re;
    _T_1843_im <= _T_1842_im;
    _T_1844_re <= _T_1843_re;
    _T_1844_im <= _T_1843_im;
    _T_1845_re <= _T_1844_re;
    _T_1845_im <= _T_1844_im;
    _T_1846_re <= _T_1845_re;
    _T_1846_im <= _T_1845_im;
    _T_1847_re <= _T_1846_re;
    _T_1847_im <= _T_1846_im;
    _T_1848_re <= _T_1847_re;
    _T_1848_im <= _T_1847_im;
    _T_1849_re <= _T_1848_re;
    _T_1849_im <= _T_1848_im;
    _T_1850_re <= _T_1849_re;
    _T_1850_im <= _T_1849_im;
    _T_1851_re <= _T_1850_re;
    _T_1851_im <= _T_1850_im;
    _T_1852_re <= _T_1851_re;
    _T_1852_im <= _T_1851_im;
    _T_1853_re <= _T_1852_re;
    _T_1853_im <= _T_1852_im;
    _T_1854_re <= _T_1853_re;
    _T_1854_im <= _T_1853_im;
    _T_1855_re <= _T_1854_re;
    _T_1855_im <= _T_1854_im;
    _T_1856_re <= _T_1855_re;
    _T_1856_im <= _T_1855_im;
    _T_1857_re <= _T_1856_re;
    _T_1857_im <= _T_1856_im;
    _T_1858_re <= _T_1857_re;
    _T_1858_im <= _T_1857_im;
    _T_1859_re <= _T_1858_re;
    _T_1859_im <= _T_1858_im;
    _T_1860_re <= _T_1859_re;
    _T_1860_im <= _T_1859_im;
    _T_1861_re <= _T_1860_re;
    _T_1861_im <= _T_1860_im;
    _T_1862_re <= _T_1861_re;
    _T_1862_im <= _T_1861_im;
    _T_1863_re <= _T_1862_re;
    _T_1863_im <= _T_1862_im;
    _T_1864_re <= _T_1863_re;
    _T_1864_im <= _T_1863_im;
    _T_1865_re <= _T_1864_re;
    _T_1865_im <= _T_1864_im;
    _T_1866_re <= _T_1865_re;
    _T_1866_im <= _T_1865_im;
    _T_1867_re <= _T_1866_re;
    _T_1867_im <= _T_1866_im;
    _T_1868_re <= _T_1867_re;
    _T_1868_im <= _T_1867_im;
    _T_1869_re <= _T_1868_re;
    _T_1869_im <= _T_1868_im;
    _T_1870_re <= _T_1869_re;
    _T_1870_im <= _T_1869_im;
    _T_1871_re <= _T_1870_re;
    _T_1871_im <= _T_1870_im;
    _T_1872_re <= _T_1871_re;
    _T_1872_im <= _T_1871_im;
    _T_1873_re <= _T_1872_re;
    _T_1873_im <= _T_1872_im;
    _T_1874_re <= _T_1873_re;
    _T_1874_im <= _T_1873_im;
    _T_1875_re <= _T_1874_re;
    _T_1875_im <= _T_1874_im;
    _T_1876_re <= _T_1875_re;
    _T_1876_im <= _T_1875_im;
    _T_1877_re <= _T_1876_re;
    _T_1877_im <= _T_1876_im;
    _T_1878_re <= _T_1877_re;
    _T_1878_im <= _T_1877_im;
    _T_1879_re <= _T_1878_re;
    _T_1879_im <= _T_1878_im;
    _T_1880_re <= _T_1879_re;
    _T_1880_im <= _T_1879_im;
    _T_1881_re <= _T_1880_re;
    _T_1881_im <= _T_1880_im;
    _T_1882_re <= _T_1881_re;
    _T_1882_im <= _T_1881_im;
    _T_1883_re <= _T_1882_re;
    _T_1883_im <= _T_1882_im;
    _T_1884_re <= _T_1883_re;
    _T_1884_im <= _T_1883_im;
    _T_1885_re <= _T_1884_re;
    _T_1885_im <= _T_1884_im;
    _T_1886_re <= _T_1885_re;
    _T_1886_im <= _T_1885_im;
    _T_1887_re <= _T_1886_re;
    _T_1887_im <= _T_1886_im;
    _T_1888_re <= _T_1887_re;
    _T_1888_im <= _T_1887_im;
    _T_1889_re <= _T_1888_re;
    _T_1889_im <= _T_1888_im;
    _T_1890_re <= _T_1889_re;
    _T_1890_im <= _T_1889_im;
    _T_1891_re <= _T_1890_re;
    _T_1891_im <= _T_1890_im;
    _T_1892_re <= _T_1891_re;
    _T_1892_im <= _T_1891_im;
    _T_1893_re <= _T_1892_re;
    _T_1893_im <= _T_1892_im;
    _T_1894_re <= _T_1893_re;
    _T_1894_im <= _T_1893_im;
    _T_1895_re <= _T_1894_re;
    _T_1895_im <= _T_1894_im;
    _T_1896_re <= _T_1895_re;
    _T_1896_im <= _T_1895_im;
    _T_1897_re <= _T_1896_re;
    _T_1897_im <= _T_1896_im;
    _T_1898_re <= _T_1897_re;
    _T_1898_im <= _T_1897_im;
    _T_1899_re <= _T_1898_re;
    _T_1899_im <= _T_1898_im;
    _T_1900_re <= _T_1899_re;
    _T_1900_im <= _T_1899_im;
    _T_1901_re <= _T_1900_re;
    _T_1901_im <= _T_1900_im;
    _T_1902_re <= _T_1901_re;
    _T_1902_im <= _T_1901_im;
    _T_1903_re <= _T_1902_re;
    _T_1903_im <= _T_1902_im;
    _T_1904_re <= _T_1903_re;
    _T_1904_im <= _T_1903_im;
    _T_1905_re <= _T_1904_re;
    _T_1905_im <= _T_1904_im;
    _T_1906_re <= _T_1905_re;
    _T_1906_im <= _T_1905_im;
    _T_1907_re <= _T_1906_re;
    _T_1907_im <= _T_1906_im;
    _T_1908_re <= _T_1907_re;
    _T_1908_im <= _T_1907_im;
    _T_1909_re <= _T_1908_re;
    _T_1909_im <= _T_1908_im;
    _T_1910_re <= _T_1909_re;
    _T_1910_im <= _T_1909_im;
    _T_1911_re <= _T_1910_re;
    _T_1911_im <= _T_1910_im;
    _T_1912_re <= _T_1911_re;
    _T_1912_im <= _T_1911_im;
    _T_1913_re <= _T_1912_re;
    _T_1913_im <= _T_1912_im;
    _T_1914_re <= _T_1913_re;
    _T_1914_im <= _T_1913_im;
    _T_1915_re <= _T_1914_re;
    _T_1915_im <= _T_1914_im;
    _T_1916_re <= _T_1915_re;
    _T_1916_im <= _T_1915_im;
    _T_1917_re <= _T_1916_re;
    _T_1917_im <= _T_1916_im;
    _T_1918_re <= _T_1917_re;
    _T_1918_im <= _T_1917_im;
    _T_1919_re <= _T_1918_re;
    _T_1919_im <= _T_1918_im;
    _T_1920_re <= _T_1919_re;
    _T_1920_im <= _T_1919_im;
    _T_1921_re <= _T_1920_re;
    _T_1921_im <= _T_1920_im;
    _T_1922_re <= _T_1921_re;
    _T_1922_im <= _T_1921_im;
    _T_1923_re <= _T_1922_re;
    _T_1923_im <= _T_1922_im;
    _T_1924_re <= _T_1923_re;
    _T_1924_im <= _T_1923_im;
    _T_1925_re <= _T_1924_re;
    _T_1925_im <= _T_1924_im;
    _T_1926_re <= _T_1925_re;
    _T_1926_im <= _T_1925_im;
    _T_1927_re <= _T_1926_re;
    _T_1927_im <= _T_1926_im;
    _T_1928_re <= _T_1927_re;
    _T_1928_im <= _T_1927_im;
    _T_1929_re <= _T_1928_re;
    _T_1929_im <= _T_1928_im;
    _T_1930_re <= _T_1929_re;
    _T_1930_im <= _T_1929_im;
    _T_1931_re <= _T_1930_re;
    _T_1931_im <= _T_1930_im;
    _T_1932_re <= _T_1931_re;
    _T_1932_im <= _T_1931_im;
    _T_1933_re <= _T_1932_re;
    _T_1933_im <= _T_1932_im;
    _T_1934_re <= _T_1933_re;
    _T_1934_im <= _T_1933_im;
    _T_1935_re <= _T_1934_re;
    _T_1935_im <= _T_1934_im;
    _T_1936_re <= _T_1935_re;
    _T_1936_im <= _T_1935_im;
    _T_1937_re <= _T_1936_re;
    _T_1937_im <= _T_1936_im;
    _T_1938_re <= _T_1937_re;
    _T_1938_im <= _T_1937_im;
    _T_1939_re <= _T_1938_re;
    _T_1939_im <= _T_1938_im;
    _T_1940_re <= _T_1939_re;
    _T_1940_im <= _T_1939_im;
    _T_1941_re <= _T_1940_re;
    _T_1941_im <= _T_1940_im;
    _T_1942_re <= _T_1941_re;
    _T_1942_im <= _T_1941_im;
    _T_1943_re <= _T_1942_re;
    _T_1943_im <= _T_1942_im;
    _T_1944_re <= _T_1943_re;
    _T_1944_im <= _T_1943_im;
    _T_1945_re <= _T_1944_re;
    _T_1945_im <= _T_1944_im;
    _T_1946_re <= _T_1945_re;
    _T_1946_im <= _T_1945_im;
    _T_1947_re <= _T_1946_re;
    _T_1947_im <= _T_1946_im;
    _T_1948_re <= _T_1947_re;
    _T_1948_im <= _T_1947_im;
    _T_1949_re <= _T_1948_re;
    _T_1949_im <= _T_1948_im;
    _T_1950_re <= _T_1949_re;
    _T_1950_im <= _T_1949_im;
    _T_1951_re <= _T_1950_re;
    _T_1951_im <= _T_1950_im;
    _T_1952_re <= _T_1951_re;
    _T_1952_im <= _T_1951_im;
    _T_1953_re <= _T_1952_re;
    _T_1953_im <= _T_1952_im;
    _T_1954_re <= _T_1953_re;
    _T_1954_im <= _T_1953_im;
    _T_1955_re <= _T_1954_re;
    _T_1955_im <= _T_1954_im;
    _T_1956_re <= _T_1955_re;
    _T_1956_im <= _T_1955_im;
    _T_1957_re <= _T_1956_re;
    _T_1957_im <= _T_1956_im;
    _T_1958_re <= _T_1957_re;
    _T_1958_im <= _T_1957_im;
    _T_1959_re <= _T_1958_re;
    _T_1959_im <= _T_1958_im;
    _T_1960_re <= _T_1959_re;
    _T_1960_im <= _T_1959_im;
    _T_1961_re <= _T_1960_re;
    _T_1961_im <= _T_1960_im;
    _T_1962_re <= _T_1961_re;
    _T_1962_im <= _T_1961_im;
    _T_1963_re <= _T_1962_re;
    _T_1963_im <= _T_1962_im;
    _T_1964_re <= _T_1963_re;
    _T_1964_im <= _T_1963_im;
    _T_1965_re <= _T_1964_re;
    _T_1965_im <= _T_1964_im;
    _T_1966_re <= _T_1965_re;
    _T_1966_im <= _T_1965_im;
    _T_1967_re <= _T_1966_re;
    _T_1967_im <= _T_1966_im;
    _T_1968_re <= _T_1967_re;
    _T_1968_im <= _T_1967_im;
    _T_1969_re <= _T_1968_re;
    _T_1969_im <= _T_1968_im;
    _T_1970_re <= _T_1969_re;
    _T_1970_im <= _T_1969_im;
    _T_1971_re <= _T_1970_re;
    _T_1971_im <= _T_1970_im;
    _T_1972_re <= _T_1971_re;
    _T_1972_im <= _T_1971_im;
    _T_1973_re <= _T_1972_re;
    _T_1973_im <= _T_1972_im;
    _T_1974_re <= _T_1973_re;
    _T_1974_im <= _T_1973_im;
    _T_1975_re <= _T_1974_re;
    _T_1975_im <= _T_1974_im;
    _T_1976_re <= _T_1975_re;
    _T_1976_im <= _T_1975_im;
    _T_1977_re <= _T_1976_re;
    _T_1977_im <= _T_1976_im;
    _T_1978_re <= _T_1977_re;
    _T_1978_im <= _T_1977_im;
    _T_1979_re <= _T_1978_re;
    _T_1979_im <= _T_1978_im;
    _T_1980_re <= _T_1979_re;
    _T_1980_im <= _T_1979_im;
    _T_1981_re <= _T_1980_re;
    _T_1981_im <= _T_1980_im;
    _T_1982_re <= _T_1981_re;
    _T_1982_im <= _T_1981_im;
    _T_1983_re <= _T_1982_re;
    _T_1983_im <= _T_1982_im;
    _T_1984_re <= _T_1983_re;
    _T_1984_im <= _T_1983_im;
    _T_1985_re <= _T_1984_re;
    _T_1985_im <= _T_1984_im;
    _T_1986_re <= _T_1985_re;
    _T_1986_im <= _T_1985_im;
    _T_1987_re <= _T_1986_re;
    _T_1987_im <= _T_1986_im;
    _T_1988_re <= _T_1987_re;
    _T_1988_im <= _T_1987_im;
    _T_1989_re <= _T_1988_re;
    _T_1989_im <= _T_1988_im;
    _T_1990_re <= _T_1989_re;
    _T_1990_im <= _T_1989_im;
    _T_1991_re <= _T_1990_re;
    _T_1991_im <= _T_1990_im;
    _T_1992_re <= _T_1991_re;
    _T_1992_im <= _T_1991_im;
    _T_1993_re <= _T_1992_re;
    _T_1993_im <= _T_1992_im;
    _T_1994_re <= _T_1993_re;
    _T_1994_im <= _T_1993_im;
    _T_1995_re <= _T_1994_re;
    _T_1995_im <= _T_1994_im;
    _T_1996_re <= _T_1995_re;
    _T_1996_im <= _T_1995_im;
    _T_1997_re <= _T_1996_re;
    _T_1997_im <= _T_1996_im;
    _T_1998_re <= _T_1997_re;
    _T_1998_im <= _T_1997_im;
    _T_1999_re <= _T_1998_re;
    _T_1999_im <= _T_1998_im;
    _T_2000_re <= _T_1999_re;
    _T_2000_im <= _T_1999_im;
    _T_2001_re <= _T_2000_re;
    _T_2001_im <= _T_2000_im;
    _T_2002_re <= _T_2001_re;
    _T_2002_im <= _T_2001_im;
    _T_2003_re <= _T_2002_re;
    _T_2003_im <= _T_2002_im;
    _T_2004_re <= _T_2003_re;
    _T_2004_im <= _T_2003_im;
    _T_2005_re <= _T_2004_re;
    _T_2005_im <= _T_2004_im;
    _T_2006_re <= _T_2005_re;
    _T_2006_im <= _T_2005_im;
    _T_2007_re <= _T_2006_re;
    _T_2007_im <= _T_2006_im;
    _T_2008_re <= _T_2007_re;
    _T_2008_im <= _T_2007_im;
    _T_2009_re <= _T_2008_re;
    _T_2009_im <= _T_2008_im;
    _T_2010_re <= _T_2009_re;
    _T_2010_im <= _T_2009_im;
    _T_2011_re <= _T_2010_re;
    _T_2011_im <= _T_2010_im;
    _T_2012_re <= _T_2011_re;
    _T_2012_im <= _T_2011_im;
    _T_2013_re <= _T_2012_re;
    _T_2013_im <= _T_2012_im;
    _T_2014_re <= _T_2013_re;
    _T_2014_im <= _T_2013_im;
    _T_2015_re <= _T_2014_re;
    _T_2015_im <= _T_2014_im;
    _T_2016_re <= _T_2015_re;
    _T_2016_im <= _T_2015_im;
    _T_2017_re <= _T_2016_re;
    _T_2017_im <= _T_2016_im;
    _T_2018_re <= _T_2017_re;
    _T_2018_im <= _T_2017_im;
    _T_2019_re <= _T_2018_re;
    _T_2019_im <= _T_2018_im;
    _T_2020_re <= _T_2019_re;
    _T_2020_im <= _T_2019_im;
    _T_2021_re <= _T_2020_re;
    _T_2021_im <= _T_2020_im;
    _T_2022_re <= _T_2021_re;
    _T_2022_im <= _T_2021_im;
    _T_2023_re <= _T_2022_re;
    _T_2023_im <= _T_2022_im;
    _T_2024_re <= _T_2023_re;
    _T_2024_im <= _T_2023_im;
    _T_2025_re <= _T_2024_re;
    _T_2025_im <= _T_2024_im;
    _T_2026_re <= _T_2025_re;
    _T_2026_im <= _T_2025_im;
    _T_2027_re <= _T_2026_re;
    _T_2027_im <= _T_2026_im;
    _T_2028_re <= _T_2027_re;
    _T_2028_im <= _T_2027_im;
    _T_2029_re <= _T_2028_re;
    _T_2029_im <= _T_2028_im;
    _T_2030_re <= _T_2029_re;
    _T_2030_im <= _T_2029_im;
    _T_2031_re <= _T_2030_re;
    _T_2031_im <= _T_2030_im;
    _T_2032_re <= _T_2031_re;
    _T_2032_im <= _T_2031_im;
    _T_2033_re <= _T_2032_re;
    _T_2033_im <= _T_2032_im;
    _T_2034_re <= _T_2033_re;
    _T_2034_im <= _T_2033_im;
    _T_2035_re <= _T_2034_re;
    _T_2035_im <= _T_2034_im;
    _T_2036_re <= _T_2035_re;
    _T_2036_im <= _T_2035_im;
    _T_2037_re <= _T_2036_re;
    _T_2037_im <= _T_2036_im;
    _T_2038_re <= _T_2037_re;
    _T_2038_im <= _T_2037_im;
    _T_2039_re <= _T_2038_re;
    _T_2039_im <= _T_2038_im;
    _T_2040_re <= _T_2039_re;
    _T_2040_im <= _T_2039_im;
    _T_2041_re <= _T_2040_re;
    _T_2041_im <= _T_2040_im;
    _T_2042_re <= _T_2041_re;
    _T_2042_im <= _T_2041_im;
    _T_2043_re <= _T_2042_re;
    _T_2043_im <= _T_2042_im;
    _T_2044_re <= _T_2043_re;
    _T_2044_im <= _T_2043_im;
    _T_2045_re <= _T_2044_re;
    _T_2045_im <= _T_2044_im;
    _T_2046_re <= _T_2045_re;
    _T_2046_im <= _T_2045_im;
    _T_2047_re <= _T_2046_re;
    _T_2047_im <= _T_2046_im;
    _T_2048_re <= _T_2047_re;
    _T_2048_im <= _T_2047_im;
    _T_2049_re <= _T_2048_re;
    _T_2049_im <= _T_2048_im;
    _T_2050_re <= _T_2049_re;
    _T_2050_im <= _T_2049_im;
    _T_2051_re <= _T_2050_re;
    _T_2051_im <= _T_2050_im;
    _T_2052_re <= _T_2051_re;
    _T_2052_im <= _T_2051_im;
    _T_2053_re <= _T_2052_re;
    _T_2053_im <= _T_2052_im;
    _T_2054_re <= _T_2053_re;
    _T_2054_im <= _T_2053_im;
    _T_2055_re <= _T_2054_re;
    _T_2055_im <= _T_2054_im;
    _T_2056_re <= _T_2055_re;
    _T_2056_im <= _T_2055_im;
    _T_2057_re <= _T_2056_re;
    _T_2057_im <= _T_2056_im;
    _T_2058_re <= _T_2057_re;
    _T_2058_im <= _T_2057_im;
    _T_2059_re <= _T_2058_re;
    _T_2059_im <= _T_2058_im;
    _T_2060_re <= _T_2059_re;
    _T_2060_im <= _T_2059_im;
    _T_2061_re <= _T_2060_re;
    _T_2061_im <= _T_2060_im;
    _T_2062_re <= _T_2061_re;
    _T_2062_im <= _T_2061_im;
    _T_2063_re <= _T_2062_re;
    _T_2063_im <= _T_2062_im;
    _T_2064_re <= _T_2063_re;
    _T_2064_im <= _T_2063_im;
    _T_2065_re <= _T_2064_re;
    _T_2065_im <= _T_2064_im;
    _T_2066_re <= _T_2065_re;
    _T_2066_im <= _T_2065_im;
    _T_2067_re <= _T_2066_re;
    _T_2067_im <= _T_2066_im;
    _T_2068_re <= _T_2067_re;
    _T_2068_im <= _T_2067_im;
    _T_2069_re <= _T_2068_re;
    _T_2069_im <= _T_2068_im;
    _T_2070_re <= _T_2069_re;
    _T_2070_im <= _T_2069_im;
    _T_2071_re <= _T_2070_re;
    _T_2071_im <= _T_2070_im;
    _T_2072_re <= _T_2071_re;
    _T_2072_im <= _T_2071_im;
    _T_2073_re <= _T_2072_re;
    _T_2073_im <= _T_2072_im;
    _T_2074_re <= _T_2073_re;
    _T_2074_im <= _T_2073_im;
    _T_2075_re <= _T_2074_re;
    _T_2075_im <= _T_2074_im;
    _T_2076_re <= _T_2075_re;
    _T_2076_im <= _T_2075_im;
    _T_2077_re <= _T_2076_re;
    _T_2077_im <= _T_2076_im;
    _T_2078_re <= _T_2077_re;
    _T_2078_im <= _T_2077_im;
    _T_2079_re <= _T_2078_re;
    _T_2079_im <= _T_2078_im;
    _T_2080_re <= _T_2079_re;
    _T_2080_im <= _T_2079_im;
    _T_2081_re <= _T_2080_re;
    _T_2081_im <= _T_2080_im;
    _T_2082_re <= _T_2081_re;
    _T_2082_im <= _T_2081_im;
    _T_2083_re <= _T_2082_re;
    _T_2083_im <= _T_2082_im;
    _T_2084_re <= _T_2083_re;
    _T_2084_im <= _T_2083_im;
    _T_2085_re <= _T_2084_re;
    _T_2085_im <= _T_2084_im;
    _T_2086_re <= _T_2085_re;
    _T_2086_im <= _T_2085_im;
    _T_2087_re <= _T_2086_re;
    _T_2087_im <= _T_2086_im;
    _T_2088_re <= _T_2087_re;
    _T_2088_im <= _T_2087_im;
    _T_2089_re <= _T_2088_re;
    _T_2089_im <= _T_2088_im;
    _T_2090_re <= _T_2089_re;
    _T_2090_im <= _T_2089_im;
    _T_2091_re <= _T_2090_re;
    _T_2091_im <= _T_2090_im;
    _T_2092_re <= _T_2091_re;
    _T_2092_im <= _T_2091_im;
    _T_2093_re <= _T_2092_re;
    _T_2093_im <= _T_2092_im;
    _T_2094_re <= _T_2093_re;
    _T_2094_im <= _T_2093_im;
    _T_2095_re <= _T_2094_re;
    _T_2095_im <= _T_2094_im;
    _T_2096_re <= _T_2095_re;
    _T_2096_im <= _T_2095_im;
    _T_2097_re <= _T_2096_re;
    _T_2097_im <= _T_2096_im;
    _T_2098_re <= _T_2097_re;
    _T_2098_im <= _T_2097_im;
    _T_2099_re <= _T_2098_re;
    _T_2099_im <= _T_2098_im;
    _T_2100_re <= _T_2099_re;
    _T_2100_im <= _T_2099_im;
    _T_2101_re <= _T_2100_re;
    _T_2101_im <= _T_2100_im;
    _T_2102_re <= _T_2101_re;
    _T_2102_im <= _T_2101_im;
    _T_2103_re <= _T_2102_re;
    _T_2103_im <= _T_2102_im;
    _T_2104_re <= _T_2103_re;
    _T_2104_im <= _T_2103_im;
    _T_2105_re <= _T_2104_re;
    _T_2105_im <= _T_2104_im;
    _T_2106_re <= _T_2105_re;
    _T_2106_im <= _T_2105_im;
    _T_2107_re <= _T_2106_re;
    _T_2107_im <= _T_2106_im;
    _T_2108_re <= _T_2107_re;
    _T_2108_im <= _T_2107_im;
    _T_2109_re <= _T_2108_re;
    _T_2109_im <= _T_2108_im;
    _T_2110_re <= _T_2109_re;
    _T_2110_im <= _T_2109_im;
    _T_2111_re <= _T_2110_re;
    _T_2111_im <= _T_2110_im;
    _T_2112_re <= _T_2111_re;
    _T_2112_im <= _T_2111_im;
    _T_2113_re <= _T_2112_re;
    _T_2113_im <= _T_2112_im;
    _T_2114_re <= _T_2113_re;
    _T_2114_im <= _T_2113_im;
    _T_2115_re <= _T_2114_re;
    _T_2115_im <= _T_2114_im;
    _T_2116_re <= _T_2115_re;
    _T_2116_im <= _T_2115_im;
    _T_2117_re <= _T_2116_re;
    _T_2117_im <= _T_2116_im;
    _T_2118_re <= _T_2117_re;
    _T_2118_im <= _T_2117_im;
    _T_2119_re <= _T_2118_re;
    _T_2119_im <= _T_2118_im;
    _T_2120_re <= _T_2119_re;
    _T_2120_im <= _T_2119_im;
    _T_2121_re <= _T_2120_re;
    _T_2121_im <= _T_2120_im;
    _T_2122_re <= _T_2121_re;
    _T_2122_im <= _T_2121_im;
    _T_2123_re <= _T_2122_re;
    _T_2123_im <= _T_2122_im;
    _T_2124_re <= _T_2123_re;
    _T_2124_im <= _T_2123_im;
    _T_2125_re <= _T_2124_re;
    _T_2125_im <= _T_2124_im;
    _T_2126_re <= _T_2125_re;
    _T_2126_im <= _T_2125_im;
    _T_2127_re <= _T_2126_re;
    _T_2127_im <= _T_2126_im;
    _T_2128_re <= _T_2127_re;
    _T_2128_im <= _T_2127_im;
    _T_2129_re <= _T_2128_re;
    _T_2129_im <= _T_2128_im;
    _T_2130_re <= _T_2129_re;
    _T_2130_im <= _T_2129_im;
    _T_2131_re <= _T_2130_re;
    _T_2131_im <= _T_2130_im;
    _T_2132_re <= _T_2131_re;
    _T_2132_im <= _T_2131_im;
    _T_2133_re <= _T_2132_re;
    _T_2133_im <= _T_2132_im;
    _T_2134_re <= _T_2133_re;
    _T_2134_im <= _T_2133_im;
    _T_2135_re <= _T_2134_re;
    _T_2135_im <= _T_2134_im;
    _T_2136_re <= _T_2135_re;
    _T_2136_im <= _T_2135_im;
    _T_2137_re <= _T_2136_re;
    _T_2137_im <= _T_2136_im;
    _T_2138_re <= _T_2137_re;
    _T_2138_im <= _T_2137_im;
    _T_2139_re <= _T_2138_re;
    _T_2139_im <= _T_2138_im;
    _T_2140_re <= _T_2139_re;
    _T_2140_im <= _T_2139_im;
    _T_2141_re <= _T_2140_re;
    _T_2141_im <= _T_2140_im;
    _T_2142_re <= _T_2141_re;
    _T_2142_im <= _T_2141_im;
    _T_2143_re <= _T_2142_re;
    _T_2143_im <= _T_2142_im;
    _T_2144_re <= _T_2143_re;
    _T_2144_im <= _T_2143_im;
    _T_2145_re <= _T_2144_re;
    _T_2145_im <= _T_2144_im;
    _T_2146_re <= _T_2145_re;
    _T_2146_im <= _T_2145_im;
    _T_2147_re <= _T_2146_re;
    _T_2147_im <= _T_2146_im;
    _T_2148_re <= _T_2147_re;
    _T_2148_im <= _T_2147_im;
    _T_2149_re <= _T_2148_re;
    _T_2149_im <= _T_2148_im;
    _T_2150_re <= _T_2149_re;
    _T_2150_im <= _T_2149_im;
    _T_2151_re <= _T_2150_re;
    _T_2151_im <= _T_2150_im;
    _T_2152_re <= _T_2151_re;
    _T_2152_im <= _T_2151_im;
    _T_2153_re <= _T_2152_re;
    _T_2153_im <= _T_2152_im;
    _T_2154_re <= _T_2153_re;
    _T_2154_im <= _T_2153_im;
    _T_2155_re <= _T_2154_re;
    _T_2155_im <= _T_2154_im;
    _T_2156_re <= _T_2155_re;
    _T_2156_im <= _T_2155_im;
    _T_2157_re <= _T_2156_re;
    _T_2157_im <= _T_2156_im;
    _T_2158_re <= _T_2157_re;
    _T_2158_im <= _T_2157_im;
    _T_2159_re <= _T_2158_re;
    _T_2159_im <= _T_2158_im;
    _T_2160_re <= _T_2159_re;
    _T_2160_im <= _T_2159_im;
    _T_2161_re <= _T_2160_re;
    _T_2161_im <= _T_2160_im;
    _T_2162_re <= _T_2161_re;
    _T_2162_im <= _T_2161_im;
    _T_2163_re <= _T_2162_re;
    _T_2163_im <= _T_2162_im;
    _T_2164_re <= _T_2163_re;
    _T_2164_im <= _T_2163_im;
    _T_2165_re <= _T_2164_re;
    _T_2165_im <= _T_2164_im;
    _T_2166_re <= _T_2165_re;
    _T_2166_im <= _T_2165_im;
    _T_2167_re <= _T_2166_re;
    _T_2167_im <= _T_2166_im;
    _T_2168_re <= _T_2167_re;
    _T_2168_im <= _T_2167_im;
    _T_2169_re <= _T_2168_re;
    _T_2169_im <= _T_2168_im;
    _T_2170_re <= _T_2169_re;
    _T_2170_im <= _T_2169_im;
    _T_2171_re <= _T_2170_re;
    _T_2171_im <= _T_2170_im;
    _T_2172_re <= _T_2171_re;
    _T_2172_im <= _T_2171_im;
    _T_2173_re <= _T_2172_re;
    _T_2173_im <= _T_2172_im;
    _T_2174_re <= _T_2173_re;
    _T_2174_im <= _T_2173_im;
    _T_2175_re <= _T_2174_re;
    _T_2175_im <= _T_2174_im;
    _T_2176_re <= _T_2175_re;
    _T_2176_im <= _T_2175_im;
    _T_2177_re <= _T_2176_re;
    _T_2177_im <= _T_2176_im;
    _T_2178_re <= _T_2177_re;
    _T_2178_im <= _T_2177_im;
    _T_2179_re <= _T_2178_re;
    _T_2179_im <= _T_2178_im;
    _T_2180_re <= _T_2179_re;
    _T_2180_im <= _T_2179_im;
    _T_2181_re <= _T_2180_re;
    _T_2181_im <= _T_2180_im;
    _T_2182_re <= _T_2181_re;
    _T_2182_im <= _T_2181_im;
    _T_2183_re <= _T_2182_re;
    _T_2183_im <= _T_2182_im;
    _T_2184_re <= _T_2183_re;
    _T_2184_im <= _T_2183_im;
    _T_2185_re <= _T_2184_re;
    _T_2185_im <= _T_2184_im;
    _T_2186_re <= _T_2185_re;
    _T_2186_im <= _T_2185_im;
    _T_2187_re <= _T_2186_re;
    _T_2187_im <= _T_2186_im;
    _T_2188_re <= _T_2187_re;
    _T_2188_im <= _T_2187_im;
    _T_2189_re <= _T_2188_re;
    _T_2189_im <= _T_2188_im;
    _T_2190_re <= _T_2189_re;
    _T_2190_im <= _T_2189_im;
    _T_2191_re <= _T_2190_re;
    _T_2191_im <= _T_2190_im;
    _T_2192_re <= _T_2191_re;
    _T_2192_im <= _T_2191_im;
    _T_2193_re <= _T_2192_re;
    _T_2193_im <= _T_2192_im;
    _T_2194_re <= _T_2193_re;
    _T_2194_im <= _T_2193_im;
    _T_2195_re <= _T_2194_re;
    _T_2195_im <= _T_2194_im;
    _T_2196_re <= _T_2195_re;
    _T_2196_im <= _T_2195_im;
    _T_2197_re <= _T_2196_re;
    _T_2197_im <= _T_2196_im;
    _T_2198_re <= _T_2197_re;
    _T_2198_im <= _T_2197_im;
    _T_2199_re <= _T_2198_re;
    _T_2199_im <= _T_2198_im;
    _T_2200_re <= _T_2199_re;
    _T_2200_im <= _T_2199_im;
    _T_2201_re <= _T_2200_re;
    _T_2201_im <= _T_2200_im;
    _T_2202_re <= _T_2201_re;
    _T_2202_im <= _T_2201_im;
    _T_2203_re <= _T_2202_re;
    _T_2203_im <= _T_2202_im;
    _T_2204_re <= _T_2203_re;
    _T_2204_im <= _T_2203_im;
    _T_2205_re <= _T_2204_re;
    _T_2205_im <= _T_2204_im;
    _T_2206_re <= _T_2205_re;
    _T_2206_im <= _T_2205_im;
    _T_2207_re <= _T_2206_re;
    _T_2207_im <= _T_2206_im;
    _T_2208_re <= _T_2207_re;
    _T_2208_im <= _T_2207_im;
    _T_2209_re <= _T_2208_re;
    _T_2209_im <= _T_2208_im;
    _T_2210_re <= _T_2209_re;
    _T_2210_im <= _T_2209_im;
    _T_2211_re <= _T_2210_re;
    _T_2211_im <= _T_2210_im;
    _T_2212_re <= _T_2211_re;
    _T_2212_im <= _T_2211_im;
    _T_2213_re <= _T_2212_re;
    _T_2213_im <= _T_2212_im;
    _T_2214_re <= _T_2213_re;
    _T_2214_im <= _T_2213_im;
    _T_2215_re <= _T_2214_re;
    _T_2215_im <= _T_2214_im;
    _T_2216_re <= _T_2215_re;
    _T_2216_im <= _T_2215_im;
    _T_2217_re <= _T_2216_re;
    _T_2217_im <= _T_2216_im;
    _T_2218_re <= _T_2217_re;
    _T_2218_im <= _T_2217_im;
    _T_2219_re <= _T_2218_re;
    _T_2219_im <= _T_2218_im;
    _T_2220_re <= _T_2219_re;
    _T_2220_im <= _T_2219_im;
    _T_2221_re <= _T_2220_re;
    _T_2221_im <= _T_2220_im;
    _T_2222_re <= _T_2221_re;
    _T_2222_im <= _T_2221_im;
    _T_2223_re <= _T_2222_re;
    _T_2223_im <= _T_2222_im;
    _T_2224_re <= _T_2223_re;
    _T_2224_im <= _T_2223_im;
    _T_2225_re <= _T_2224_re;
    _T_2225_im <= _T_2224_im;
    _T_2226_re <= _T_2225_re;
    _T_2226_im <= _T_2225_im;
    _T_2227_re <= _T_2226_re;
    _T_2227_im <= _T_2226_im;
    _T_2228_re <= _T_2227_re;
    _T_2228_im <= _T_2227_im;
    _T_2229_re <= _T_2228_re;
    _T_2229_im <= _T_2228_im;
    _T_2230_re <= _T_2229_re;
    _T_2230_im <= _T_2229_im;
    _T_2231_re <= _T_2230_re;
    _T_2231_im <= _T_2230_im;
    _T_2232_re <= _T_2231_re;
    _T_2232_im <= _T_2231_im;
    _T_2233_re <= _T_2232_re;
    _T_2233_im <= _T_2232_im;
    _T_2234_re <= _T_2233_re;
    _T_2234_im <= _T_2233_im;
    _T_2235_re <= _T_2234_re;
    _T_2235_im <= _T_2234_im;
    _T_2236_re <= _T_2235_re;
    _T_2236_im <= _T_2235_im;
    _T_2237_re <= _T_2236_re;
    _T_2237_im <= _T_2236_im;
    _T_2238_re <= _T_2237_re;
    _T_2238_im <= _T_2237_im;
    _T_2239_re <= _T_2238_re;
    _T_2239_im <= _T_2238_im;
    _T_2242_re <= Butterfly_1_io_out2_re;
    _T_2242_im <= Butterfly_1_io_out2_im;
    _T_2243_re <= _T_2242_re;
    _T_2243_im <= _T_2242_im;
    _T_2244_re <= _T_2243_re;
    _T_2244_im <= _T_2243_im;
    _T_2245_re <= _T_2244_re;
    _T_2245_im <= _T_2244_im;
    _T_2246_re <= _T_2245_re;
    _T_2246_im <= _T_2245_im;
    _T_2247_re <= _T_2246_re;
    _T_2247_im <= _T_2246_im;
    _T_2248_re <= _T_2247_re;
    _T_2248_im <= _T_2247_im;
    _T_2249_re <= _T_2248_re;
    _T_2249_im <= _T_2248_im;
    _T_2250_re <= _T_2249_re;
    _T_2250_im <= _T_2249_im;
    _T_2251_re <= _T_2250_re;
    _T_2251_im <= _T_2250_im;
    _T_2252_re <= _T_2251_re;
    _T_2252_im <= _T_2251_im;
    _T_2253_re <= _T_2252_re;
    _T_2253_im <= _T_2252_im;
    _T_2254_re <= _T_2253_re;
    _T_2254_im <= _T_2253_im;
    _T_2255_re <= _T_2254_re;
    _T_2255_im <= _T_2254_im;
    _T_2256_re <= _T_2255_re;
    _T_2256_im <= _T_2255_im;
    _T_2257_re <= _T_2256_re;
    _T_2257_im <= _T_2256_im;
    _T_2258_re <= _T_2257_re;
    _T_2258_im <= _T_2257_im;
    _T_2259_re <= _T_2258_re;
    _T_2259_im <= _T_2258_im;
    _T_2260_re <= _T_2259_re;
    _T_2260_im <= _T_2259_im;
    _T_2261_re <= _T_2260_re;
    _T_2261_im <= _T_2260_im;
    _T_2262_re <= _T_2261_re;
    _T_2262_im <= _T_2261_im;
    _T_2263_re <= _T_2262_re;
    _T_2263_im <= _T_2262_im;
    _T_2264_re <= _T_2263_re;
    _T_2264_im <= _T_2263_im;
    _T_2265_re <= _T_2264_re;
    _T_2265_im <= _T_2264_im;
    _T_2266_re <= _T_2265_re;
    _T_2266_im <= _T_2265_im;
    _T_2267_re <= _T_2266_re;
    _T_2267_im <= _T_2266_im;
    _T_2268_re <= _T_2267_re;
    _T_2268_im <= _T_2267_im;
    _T_2269_re <= _T_2268_re;
    _T_2269_im <= _T_2268_im;
    _T_2270_re <= _T_2269_re;
    _T_2270_im <= _T_2269_im;
    _T_2271_re <= _T_2270_re;
    _T_2271_im <= _T_2270_im;
    _T_2272_re <= _T_2271_re;
    _T_2272_im <= _T_2271_im;
    _T_2273_re <= _T_2272_re;
    _T_2273_im <= _T_2272_im;
    _T_2274_re <= _T_2273_re;
    _T_2274_im <= _T_2273_im;
    _T_2275_re <= _T_2274_re;
    _T_2275_im <= _T_2274_im;
    _T_2276_re <= _T_2275_re;
    _T_2276_im <= _T_2275_im;
    _T_2277_re <= _T_2276_re;
    _T_2277_im <= _T_2276_im;
    _T_2278_re <= _T_2277_re;
    _T_2278_im <= _T_2277_im;
    _T_2279_re <= _T_2278_re;
    _T_2279_im <= _T_2278_im;
    _T_2280_re <= _T_2279_re;
    _T_2280_im <= _T_2279_im;
    _T_2281_re <= _T_2280_re;
    _T_2281_im <= _T_2280_im;
    _T_2282_re <= _T_2281_re;
    _T_2282_im <= _T_2281_im;
    _T_2283_re <= _T_2282_re;
    _T_2283_im <= _T_2282_im;
    _T_2284_re <= _T_2283_re;
    _T_2284_im <= _T_2283_im;
    _T_2285_re <= _T_2284_re;
    _T_2285_im <= _T_2284_im;
    _T_2286_re <= _T_2285_re;
    _T_2286_im <= _T_2285_im;
    _T_2287_re <= _T_2286_re;
    _T_2287_im <= _T_2286_im;
    _T_2288_re <= _T_2287_re;
    _T_2288_im <= _T_2287_im;
    _T_2289_re <= _T_2288_re;
    _T_2289_im <= _T_2288_im;
    _T_2290_re <= _T_2289_re;
    _T_2290_im <= _T_2289_im;
    _T_2291_re <= _T_2290_re;
    _T_2291_im <= _T_2290_im;
    _T_2292_re <= _T_2291_re;
    _T_2292_im <= _T_2291_im;
    _T_2293_re <= _T_2292_re;
    _T_2293_im <= _T_2292_im;
    _T_2294_re <= _T_2293_re;
    _T_2294_im <= _T_2293_im;
    _T_2295_re <= _T_2294_re;
    _T_2295_im <= _T_2294_im;
    _T_2296_re <= _T_2295_re;
    _T_2296_im <= _T_2295_im;
    _T_2297_re <= _T_2296_re;
    _T_2297_im <= _T_2296_im;
    _T_2298_re <= _T_2297_re;
    _T_2298_im <= _T_2297_im;
    _T_2299_re <= _T_2298_re;
    _T_2299_im <= _T_2298_im;
    _T_2300_re <= _T_2299_re;
    _T_2300_im <= _T_2299_im;
    _T_2301_re <= _T_2300_re;
    _T_2301_im <= _T_2300_im;
    _T_2302_re <= _T_2301_re;
    _T_2302_im <= _T_2301_im;
    _T_2303_re <= _T_2302_re;
    _T_2303_im <= _T_2302_im;
    _T_2304_re <= _T_2303_re;
    _T_2304_im <= _T_2303_im;
    _T_2305_re <= _T_2304_re;
    _T_2305_im <= _T_2304_im;
    _T_2306_re <= _T_2305_re;
    _T_2306_im <= _T_2305_im;
    _T_2307_re <= _T_2306_re;
    _T_2307_im <= _T_2306_im;
    _T_2308_re <= _T_2307_re;
    _T_2308_im <= _T_2307_im;
    _T_2309_re <= _T_2308_re;
    _T_2309_im <= _T_2308_im;
    _T_2310_re <= _T_2309_re;
    _T_2310_im <= _T_2309_im;
    _T_2311_re <= _T_2310_re;
    _T_2311_im <= _T_2310_im;
    _T_2312_re <= _T_2311_re;
    _T_2312_im <= _T_2311_im;
    _T_2313_re <= _T_2312_re;
    _T_2313_im <= _T_2312_im;
    _T_2314_re <= _T_2313_re;
    _T_2314_im <= _T_2313_im;
    _T_2315_re <= _T_2314_re;
    _T_2315_im <= _T_2314_im;
    _T_2316_re <= _T_2315_re;
    _T_2316_im <= _T_2315_im;
    _T_2317_re <= _T_2316_re;
    _T_2317_im <= _T_2316_im;
    _T_2318_re <= _T_2317_re;
    _T_2318_im <= _T_2317_im;
    _T_2319_re <= _T_2318_re;
    _T_2319_im <= _T_2318_im;
    _T_2320_re <= _T_2319_re;
    _T_2320_im <= _T_2319_im;
    _T_2321_re <= _T_2320_re;
    _T_2321_im <= _T_2320_im;
    _T_2322_re <= _T_2321_re;
    _T_2322_im <= _T_2321_im;
    _T_2323_re <= _T_2322_re;
    _T_2323_im <= _T_2322_im;
    _T_2324_re <= _T_2323_re;
    _T_2324_im <= _T_2323_im;
    _T_2325_re <= _T_2324_re;
    _T_2325_im <= _T_2324_im;
    _T_2326_re <= _T_2325_re;
    _T_2326_im <= _T_2325_im;
    _T_2327_re <= _T_2326_re;
    _T_2327_im <= _T_2326_im;
    _T_2328_re <= _T_2327_re;
    _T_2328_im <= _T_2327_im;
    _T_2329_re <= _T_2328_re;
    _T_2329_im <= _T_2328_im;
    _T_2330_re <= _T_2329_re;
    _T_2330_im <= _T_2329_im;
    _T_2331_re <= _T_2330_re;
    _T_2331_im <= _T_2330_im;
    _T_2332_re <= _T_2331_re;
    _T_2332_im <= _T_2331_im;
    _T_2333_re <= _T_2332_re;
    _T_2333_im <= _T_2332_im;
    _T_2334_re <= _T_2333_re;
    _T_2334_im <= _T_2333_im;
    _T_2335_re <= _T_2334_re;
    _T_2335_im <= _T_2334_im;
    _T_2336_re <= _T_2335_re;
    _T_2336_im <= _T_2335_im;
    _T_2337_re <= _T_2336_re;
    _T_2337_im <= _T_2336_im;
    _T_2338_re <= _T_2337_re;
    _T_2338_im <= _T_2337_im;
    _T_2339_re <= _T_2338_re;
    _T_2339_im <= _T_2338_im;
    _T_2340_re <= _T_2339_re;
    _T_2340_im <= _T_2339_im;
    _T_2341_re <= _T_2340_re;
    _T_2341_im <= _T_2340_im;
    _T_2342_re <= _T_2341_re;
    _T_2342_im <= _T_2341_im;
    _T_2343_re <= _T_2342_re;
    _T_2343_im <= _T_2342_im;
    _T_2344_re <= _T_2343_re;
    _T_2344_im <= _T_2343_im;
    _T_2345_re <= _T_2344_re;
    _T_2345_im <= _T_2344_im;
    _T_2346_re <= _T_2345_re;
    _T_2346_im <= _T_2345_im;
    _T_2347_re <= _T_2346_re;
    _T_2347_im <= _T_2346_im;
    _T_2348_re <= _T_2347_re;
    _T_2348_im <= _T_2347_im;
    _T_2349_re <= _T_2348_re;
    _T_2349_im <= _T_2348_im;
    _T_2350_re <= _T_2349_re;
    _T_2350_im <= _T_2349_im;
    _T_2351_re <= _T_2350_re;
    _T_2351_im <= _T_2350_im;
    _T_2352_re <= _T_2351_re;
    _T_2352_im <= _T_2351_im;
    _T_2353_re <= _T_2352_re;
    _T_2353_im <= _T_2352_im;
    _T_2354_re <= _T_2353_re;
    _T_2354_im <= _T_2353_im;
    _T_2355_re <= _T_2354_re;
    _T_2355_im <= _T_2354_im;
    _T_2356_re <= _T_2355_re;
    _T_2356_im <= _T_2355_im;
    _T_2357_re <= _T_2356_re;
    _T_2357_im <= _T_2356_im;
    _T_2358_re <= _T_2357_re;
    _T_2358_im <= _T_2357_im;
    _T_2359_re <= _T_2358_re;
    _T_2359_im <= _T_2358_im;
    _T_2360_re <= _T_2359_re;
    _T_2360_im <= _T_2359_im;
    _T_2361_re <= _T_2360_re;
    _T_2361_im <= _T_2360_im;
    _T_2362_re <= _T_2361_re;
    _T_2362_im <= _T_2361_im;
    _T_2363_re <= _T_2362_re;
    _T_2363_im <= _T_2362_im;
    _T_2364_re <= _T_2363_re;
    _T_2364_im <= _T_2363_im;
    _T_2365_re <= _T_2364_re;
    _T_2365_im <= _T_2364_im;
    _T_2366_re <= _T_2365_re;
    _T_2366_im <= _T_2365_im;
    _T_2367_re <= _T_2366_re;
    _T_2367_im <= _T_2366_im;
    _T_2368_re <= _T_2367_re;
    _T_2368_im <= _T_2367_im;
    _T_2369_re <= _T_2368_re;
    _T_2369_im <= _T_2368_im;
    _T_2370_re <= _T_2369_re;
    _T_2370_im <= _T_2369_im;
    _T_2371_re <= _T_2370_re;
    _T_2371_im <= _T_2370_im;
    _T_2372_re <= _T_2371_re;
    _T_2372_im <= _T_2371_im;
    _T_2373_re <= _T_2372_re;
    _T_2373_im <= _T_2372_im;
    _T_2374_re <= _T_2373_re;
    _T_2374_im <= _T_2373_im;
    _T_2375_re <= _T_2374_re;
    _T_2375_im <= _T_2374_im;
    _T_2376_re <= _T_2375_re;
    _T_2376_im <= _T_2375_im;
    _T_2377_re <= _T_2376_re;
    _T_2377_im <= _T_2376_im;
    _T_2378_re <= _T_2377_re;
    _T_2378_im <= _T_2377_im;
    _T_2379_re <= _T_2378_re;
    _T_2379_im <= _T_2378_im;
    _T_2380_re <= _T_2379_re;
    _T_2380_im <= _T_2379_im;
    _T_2381_re <= _T_2380_re;
    _T_2381_im <= _T_2380_im;
    _T_2382_re <= _T_2381_re;
    _T_2382_im <= _T_2381_im;
    _T_2383_re <= _T_2382_re;
    _T_2383_im <= _T_2382_im;
    _T_2384_re <= _T_2383_re;
    _T_2384_im <= _T_2383_im;
    _T_2385_re <= _T_2384_re;
    _T_2385_im <= _T_2384_im;
    _T_2386_re <= _T_2385_re;
    _T_2386_im <= _T_2385_im;
    _T_2387_re <= _T_2386_re;
    _T_2387_im <= _T_2386_im;
    _T_2388_re <= _T_2387_re;
    _T_2388_im <= _T_2387_im;
    _T_2389_re <= _T_2388_re;
    _T_2389_im <= _T_2388_im;
    _T_2390_re <= _T_2389_re;
    _T_2390_im <= _T_2389_im;
    _T_2391_re <= _T_2390_re;
    _T_2391_im <= _T_2390_im;
    _T_2392_re <= _T_2391_re;
    _T_2392_im <= _T_2391_im;
    _T_2393_re <= _T_2392_re;
    _T_2393_im <= _T_2392_im;
    _T_2394_re <= _T_2393_re;
    _T_2394_im <= _T_2393_im;
    _T_2395_re <= _T_2394_re;
    _T_2395_im <= _T_2394_im;
    _T_2396_re <= _T_2395_re;
    _T_2396_im <= _T_2395_im;
    _T_2397_re <= _T_2396_re;
    _T_2397_im <= _T_2396_im;
    _T_2398_re <= _T_2397_re;
    _T_2398_im <= _T_2397_im;
    _T_2399_re <= _T_2398_re;
    _T_2399_im <= _T_2398_im;
    _T_2400_re <= _T_2399_re;
    _T_2400_im <= _T_2399_im;
    _T_2401_re <= _T_2400_re;
    _T_2401_im <= _T_2400_im;
    _T_2402_re <= _T_2401_re;
    _T_2402_im <= _T_2401_im;
    _T_2403_re <= _T_2402_re;
    _T_2403_im <= _T_2402_im;
    _T_2404_re <= _T_2403_re;
    _T_2404_im <= _T_2403_im;
    _T_2405_re <= _T_2404_re;
    _T_2405_im <= _T_2404_im;
    _T_2406_re <= _T_2405_re;
    _T_2406_im <= _T_2405_im;
    _T_2407_re <= _T_2406_re;
    _T_2407_im <= _T_2406_im;
    _T_2408_re <= _T_2407_re;
    _T_2408_im <= _T_2407_im;
    _T_2409_re <= _T_2408_re;
    _T_2409_im <= _T_2408_im;
    _T_2410_re <= _T_2409_re;
    _T_2410_im <= _T_2409_im;
    _T_2411_re <= _T_2410_re;
    _T_2411_im <= _T_2410_im;
    _T_2412_re <= _T_2411_re;
    _T_2412_im <= _T_2411_im;
    _T_2413_re <= _T_2412_re;
    _T_2413_im <= _T_2412_im;
    _T_2414_re <= _T_2413_re;
    _T_2414_im <= _T_2413_im;
    _T_2415_re <= _T_2414_re;
    _T_2415_im <= _T_2414_im;
    _T_2416_re <= _T_2415_re;
    _T_2416_im <= _T_2415_im;
    _T_2417_re <= _T_2416_re;
    _T_2417_im <= _T_2416_im;
    _T_2418_re <= _T_2417_re;
    _T_2418_im <= _T_2417_im;
    _T_2419_re <= _T_2418_re;
    _T_2419_im <= _T_2418_im;
    _T_2420_re <= _T_2419_re;
    _T_2420_im <= _T_2419_im;
    _T_2421_re <= _T_2420_re;
    _T_2421_im <= _T_2420_im;
    _T_2422_re <= _T_2421_re;
    _T_2422_im <= _T_2421_im;
    _T_2423_re <= _T_2422_re;
    _T_2423_im <= _T_2422_im;
    _T_2424_re <= _T_2423_re;
    _T_2424_im <= _T_2423_im;
    _T_2425_re <= _T_2424_re;
    _T_2425_im <= _T_2424_im;
    _T_2426_re <= _T_2425_re;
    _T_2426_im <= _T_2425_im;
    _T_2427_re <= _T_2426_re;
    _T_2427_im <= _T_2426_im;
    _T_2428_re <= _T_2427_re;
    _T_2428_im <= _T_2427_im;
    _T_2429_re <= _T_2428_re;
    _T_2429_im <= _T_2428_im;
    _T_2430_re <= _T_2429_re;
    _T_2430_im <= _T_2429_im;
    _T_2431_re <= _T_2430_re;
    _T_2431_im <= _T_2430_im;
    _T_2432_re <= _T_2431_re;
    _T_2432_im <= _T_2431_im;
    _T_2433_re <= _T_2432_re;
    _T_2433_im <= _T_2432_im;
    _T_2434_re <= _T_2433_re;
    _T_2434_im <= _T_2433_im;
    _T_2435_re <= _T_2434_re;
    _T_2435_im <= _T_2434_im;
    _T_2436_re <= _T_2435_re;
    _T_2436_im <= _T_2435_im;
    _T_2437_re <= _T_2436_re;
    _T_2437_im <= _T_2436_im;
    _T_2438_re <= _T_2437_re;
    _T_2438_im <= _T_2437_im;
    _T_2439_re <= _T_2438_re;
    _T_2439_im <= _T_2438_im;
    _T_2440_re <= _T_2439_re;
    _T_2440_im <= _T_2439_im;
    _T_2441_re <= _T_2440_re;
    _T_2441_im <= _T_2440_im;
    _T_2442_re <= _T_2441_re;
    _T_2442_im <= _T_2441_im;
    _T_2443_re <= _T_2442_re;
    _T_2443_im <= _T_2442_im;
    _T_2444_re <= _T_2443_re;
    _T_2444_im <= _T_2443_im;
    _T_2445_re <= _T_2444_re;
    _T_2445_im <= _T_2444_im;
    _T_2446_re <= _T_2445_re;
    _T_2446_im <= _T_2445_im;
    _T_2447_re <= _T_2446_re;
    _T_2447_im <= _T_2446_im;
    _T_2448_re <= _T_2447_re;
    _T_2448_im <= _T_2447_im;
    _T_2449_re <= _T_2448_re;
    _T_2449_im <= _T_2448_im;
    _T_2450_re <= _T_2449_re;
    _T_2450_im <= _T_2449_im;
    _T_2451_re <= _T_2450_re;
    _T_2451_im <= _T_2450_im;
    _T_2452_re <= _T_2451_re;
    _T_2452_im <= _T_2451_im;
    _T_2453_re <= _T_2452_re;
    _T_2453_im <= _T_2452_im;
    _T_2454_re <= _T_2453_re;
    _T_2454_im <= _T_2453_im;
    _T_2455_re <= _T_2454_re;
    _T_2455_im <= _T_2454_im;
    _T_2456_re <= _T_2455_re;
    _T_2456_im <= _T_2455_im;
    _T_2457_re <= _T_2456_re;
    _T_2457_im <= _T_2456_im;
    _T_2458_re <= _T_2457_re;
    _T_2458_im <= _T_2457_im;
    _T_2459_re <= _T_2458_re;
    _T_2459_im <= _T_2458_im;
    _T_2460_re <= _T_2459_re;
    _T_2460_im <= _T_2459_im;
    _T_2461_re <= _T_2460_re;
    _T_2461_im <= _T_2460_im;
    _T_2462_re <= _T_2461_re;
    _T_2462_im <= _T_2461_im;
    _T_2463_re <= _T_2462_re;
    _T_2463_im <= _T_2462_im;
    _T_2464_re <= _T_2463_re;
    _T_2464_im <= _T_2463_im;
    _T_2465_re <= _T_2464_re;
    _T_2465_im <= _T_2464_im;
    _T_2466_re <= _T_2465_re;
    _T_2466_im <= _T_2465_im;
    _T_2467_re <= _T_2466_re;
    _T_2467_im <= _T_2466_im;
    _T_2468_re <= _T_2467_re;
    _T_2468_im <= _T_2467_im;
    _T_2469_re <= _T_2468_re;
    _T_2469_im <= _T_2468_im;
    _T_2470_re <= _T_2469_re;
    _T_2470_im <= _T_2469_im;
    _T_2471_re <= _T_2470_re;
    _T_2471_im <= _T_2470_im;
    _T_2472_re <= _T_2471_re;
    _T_2472_im <= _T_2471_im;
    _T_2473_re <= _T_2472_re;
    _T_2473_im <= _T_2472_im;
    _T_2474_re <= _T_2473_re;
    _T_2474_im <= _T_2473_im;
    _T_2475_re <= _T_2474_re;
    _T_2475_im <= _T_2474_im;
    _T_2476_re <= _T_2475_re;
    _T_2476_im <= _T_2475_im;
    _T_2477_re <= _T_2476_re;
    _T_2477_im <= _T_2476_im;
    _T_2478_re <= _T_2477_re;
    _T_2478_im <= _T_2477_im;
    _T_2479_re <= _T_2478_re;
    _T_2479_im <= _T_2478_im;
    _T_2480_re <= _T_2479_re;
    _T_2480_im <= _T_2479_im;
    _T_2481_re <= _T_2480_re;
    _T_2481_im <= _T_2480_im;
    _T_2482_re <= _T_2481_re;
    _T_2482_im <= _T_2481_im;
    _T_2483_re <= _T_2482_re;
    _T_2483_im <= _T_2482_im;
    _T_2484_re <= _T_2483_re;
    _T_2484_im <= _T_2483_im;
    _T_2485_re <= _T_2484_re;
    _T_2485_im <= _T_2484_im;
    _T_2486_re <= _T_2485_re;
    _T_2486_im <= _T_2485_im;
    _T_2487_re <= _T_2486_re;
    _T_2487_im <= _T_2486_im;
    _T_2488_re <= _T_2487_re;
    _T_2488_im <= _T_2487_im;
    _T_2489_re <= _T_2488_re;
    _T_2489_im <= _T_2488_im;
    _T_2490_re <= _T_2489_re;
    _T_2490_im <= _T_2489_im;
    _T_2491_re <= _T_2490_re;
    _T_2491_im <= _T_2490_im;
    _T_2492_re <= _T_2491_re;
    _T_2492_im <= _T_2491_im;
    _T_2493_re <= _T_2492_re;
    _T_2493_im <= _T_2492_im;
    _T_2494_re <= _T_2493_re;
    _T_2494_im <= _T_2493_im;
    _T_2495_re <= _T_2494_re;
    _T_2495_im <= _T_2494_im;
    _T_2496_re <= _T_2495_re;
    _T_2496_im <= _T_2495_im;
    _T_2497_re <= _T_2496_re;
    _T_2497_im <= _T_2496_im;
    _T_2507_re <= Switch_1_io_out1_re;
    _T_2507_im <= Switch_1_io_out1_im;
    _T_2508_re <= _T_2507_re;
    _T_2508_im <= _T_2507_im;
    _T_2509_re <= _T_2508_re;
    _T_2509_im <= _T_2508_im;
    _T_2510_re <= _T_2509_re;
    _T_2510_im <= _T_2509_im;
    _T_2511_re <= _T_2510_re;
    _T_2511_im <= _T_2510_im;
    _T_2512_re <= _T_2511_re;
    _T_2512_im <= _T_2511_im;
    _T_2513_re <= _T_2512_re;
    _T_2513_im <= _T_2512_im;
    _T_2514_re <= _T_2513_re;
    _T_2514_im <= _T_2513_im;
    _T_2515_re <= _T_2514_re;
    _T_2515_im <= _T_2514_im;
    _T_2516_re <= _T_2515_re;
    _T_2516_im <= _T_2515_im;
    _T_2517_re <= _T_2516_re;
    _T_2517_im <= _T_2516_im;
    _T_2518_re <= _T_2517_re;
    _T_2518_im <= _T_2517_im;
    _T_2519_re <= _T_2518_re;
    _T_2519_im <= _T_2518_im;
    _T_2520_re <= _T_2519_re;
    _T_2520_im <= _T_2519_im;
    _T_2521_re <= _T_2520_re;
    _T_2521_im <= _T_2520_im;
    _T_2522_re <= _T_2521_re;
    _T_2522_im <= _T_2521_im;
    _T_2523_re <= _T_2522_re;
    _T_2523_im <= _T_2522_im;
    _T_2524_re <= _T_2523_re;
    _T_2524_im <= _T_2523_im;
    _T_2525_re <= _T_2524_re;
    _T_2525_im <= _T_2524_im;
    _T_2526_re <= _T_2525_re;
    _T_2526_im <= _T_2525_im;
    _T_2527_re <= _T_2526_re;
    _T_2527_im <= _T_2526_im;
    _T_2528_re <= _T_2527_re;
    _T_2528_im <= _T_2527_im;
    _T_2529_re <= _T_2528_re;
    _T_2529_im <= _T_2528_im;
    _T_2530_re <= _T_2529_re;
    _T_2530_im <= _T_2529_im;
    _T_2531_re <= _T_2530_re;
    _T_2531_im <= _T_2530_im;
    _T_2532_re <= _T_2531_re;
    _T_2532_im <= _T_2531_im;
    _T_2533_re <= _T_2532_re;
    _T_2533_im <= _T_2532_im;
    _T_2534_re <= _T_2533_re;
    _T_2534_im <= _T_2533_im;
    _T_2535_re <= _T_2534_re;
    _T_2535_im <= _T_2534_im;
    _T_2536_re <= _T_2535_re;
    _T_2536_im <= _T_2535_im;
    _T_2537_re <= _T_2536_re;
    _T_2537_im <= _T_2536_im;
    _T_2538_re <= _T_2537_re;
    _T_2538_im <= _T_2537_im;
    _T_2539_re <= _T_2538_re;
    _T_2539_im <= _T_2538_im;
    _T_2540_re <= _T_2539_re;
    _T_2540_im <= _T_2539_im;
    _T_2541_re <= _T_2540_re;
    _T_2541_im <= _T_2540_im;
    _T_2542_re <= _T_2541_re;
    _T_2542_im <= _T_2541_im;
    _T_2543_re <= _T_2542_re;
    _T_2543_im <= _T_2542_im;
    _T_2544_re <= _T_2543_re;
    _T_2544_im <= _T_2543_im;
    _T_2545_re <= _T_2544_re;
    _T_2545_im <= _T_2544_im;
    _T_2546_re <= _T_2545_re;
    _T_2546_im <= _T_2545_im;
    _T_2547_re <= _T_2546_re;
    _T_2547_im <= _T_2546_im;
    _T_2548_re <= _T_2547_re;
    _T_2548_im <= _T_2547_im;
    _T_2549_re <= _T_2548_re;
    _T_2549_im <= _T_2548_im;
    _T_2550_re <= _T_2549_re;
    _T_2550_im <= _T_2549_im;
    _T_2551_re <= _T_2550_re;
    _T_2551_im <= _T_2550_im;
    _T_2552_re <= _T_2551_re;
    _T_2552_im <= _T_2551_im;
    _T_2553_re <= _T_2552_re;
    _T_2553_im <= _T_2552_im;
    _T_2554_re <= _T_2553_re;
    _T_2554_im <= _T_2553_im;
    _T_2555_re <= _T_2554_re;
    _T_2555_im <= _T_2554_im;
    _T_2556_re <= _T_2555_re;
    _T_2556_im <= _T_2555_im;
    _T_2557_re <= _T_2556_re;
    _T_2557_im <= _T_2556_im;
    _T_2558_re <= _T_2557_re;
    _T_2558_im <= _T_2557_im;
    _T_2559_re <= _T_2558_re;
    _T_2559_im <= _T_2558_im;
    _T_2560_re <= _T_2559_re;
    _T_2560_im <= _T_2559_im;
    _T_2561_re <= _T_2560_re;
    _T_2561_im <= _T_2560_im;
    _T_2562_re <= _T_2561_re;
    _T_2562_im <= _T_2561_im;
    _T_2563_re <= _T_2562_re;
    _T_2563_im <= _T_2562_im;
    _T_2564_re <= _T_2563_re;
    _T_2564_im <= _T_2563_im;
    _T_2565_re <= _T_2564_re;
    _T_2565_im <= _T_2564_im;
    _T_2566_re <= _T_2565_re;
    _T_2566_im <= _T_2565_im;
    _T_2567_re <= _T_2566_re;
    _T_2567_im <= _T_2566_im;
    _T_2568_re <= _T_2567_re;
    _T_2568_im <= _T_2567_im;
    _T_2569_re <= _T_2568_re;
    _T_2569_im <= _T_2568_im;
    _T_2570_re <= _T_2569_re;
    _T_2570_im <= _T_2569_im;
    _T_2571_re <= _T_2570_re;
    _T_2571_im <= _T_2570_im;
    _T_2572_re <= _T_2571_re;
    _T_2572_im <= _T_2571_im;
    _T_2573_re <= _T_2572_re;
    _T_2573_im <= _T_2572_im;
    _T_2574_re <= _T_2573_re;
    _T_2574_im <= _T_2573_im;
    _T_2575_re <= _T_2574_re;
    _T_2575_im <= _T_2574_im;
    _T_2576_re <= _T_2575_re;
    _T_2576_im <= _T_2575_im;
    _T_2577_re <= _T_2576_re;
    _T_2577_im <= _T_2576_im;
    _T_2578_re <= _T_2577_re;
    _T_2578_im <= _T_2577_im;
    _T_2579_re <= _T_2578_re;
    _T_2579_im <= _T_2578_im;
    _T_2580_re <= _T_2579_re;
    _T_2580_im <= _T_2579_im;
    _T_2581_re <= _T_2580_re;
    _T_2581_im <= _T_2580_im;
    _T_2582_re <= _T_2581_re;
    _T_2582_im <= _T_2581_im;
    _T_2583_re <= _T_2582_re;
    _T_2583_im <= _T_2582_im;
    _T_2584_re <= _T_2583_re;
    _T_2584_im <= _T_2583_im;
    _T_2585_re <= _T_2584_re;
    _T_2585_im <= _T_2584_im;
    _T_2586_re <= _T_2585_re;
    _T_2586_im <= _T_2585_im;
    _T_2587_re <= _T_2586_re;
    _T_2587_im <= _T_2586_im;
    _T_2588_re <= _T_2587_re;
    _T_2588_im <= _T_2587_im;
    _T_2589_re <= _T_2588_re;
    _T_2589_im <= _T_2588_im;
    _T_2590_re <= _T_2589_re;
    _T_2590_im <= _T_2589_im;
    _T_2591_re <= _T_2590_re;
    _T_2591_im <= _T_2590_im;
    _T_2592_re <= _T_2591_re;
    _T_2592_im <= _T_2591_im;
    _T_2593_re <= _T_2592_re;
    _T_2593_im <= _T_2592_im;
    _T_2594_re <= _T_2593_re;
    _T_2594_im <= _T_2593_im;
    _T_2595_re <= _T_2594_re;
    _T_2595_im <= _T_2594_im;
    _T_2596_re <= _T_2595_re;
    _T_2596_im <= _T_2595_im;
    _T_2597_re <= _T_2596_re;
    _T_2597_im <= _T_2596_im;
    _T_2598_re <= _T_2597_re;
    _T_2598_im <= _T_2597_im;
    _T_2599_re <= _T_2598_re;
    _T_2599_im <= _T_2598_im;
    _T_2600_re <= _T_2599_re;
    _T_2600_im <= _T_2599_im;
    _T_2601_re <= _T_2600_re;
    _T_2601_im <= _T_2600_im;
    _T_2602_re <= _T_2601_re;
    _T_2602_im <= _T_2601_im;
    _T_2603_re <= _T_2602_re;
    _T_2603_im <= _T_2602_im;
    _T_2604_re <= _T_2603_re;
    _T_2604_im <= _T_2603_im;
    _T_2605_re <= _T_2604_re;
    _T_2605_im <= _T_2604_im;
    _T_2606_re <= _T_2605_re;
    _T_2606_im <= _T_2605_im;
    _T_2607_re <= _T_2606_re;
    _T_2607_im <= _T_2606_im;
    _T_2608_re <= _T_2607_re;
    _T_2608_im <= _T_2607_im;
    _T_2609_re <= _T_2608_re;
    _T_2609_im <= _T_2608_im;
    _T_2610_re <= _T_2609_re;
    _T_2610_im <= _T_2609_im;
    _T_2611_re <= _T_2610_re;
    _T_2611_im <= _T_2610_im;
    _T_2612_re <= _T_2611_re;
    _T_2612_im <= _T_2611_im;
    _T_2613_re <= _T_2612_re;
    _T_2613_im <= _T_2612_im;
    _T_2614_re <= _T_2613_re;
    _T_2614_im <= _T_2613_im;
    _T_2615_re <= _T_2614_re;
    _T_2615_im <= _T_2614_im;
    _T_2616_re <= _T_2615_re;
    _T_2616_im <= _T_2615_im;
    _T_2617_re <= _T_2616_re;
    _T_2617_im <= _T_2616_im;
    _T_2618_re <= _T_2617_re;
    _T_2618_im <= _T_2617_im;
    _T_2619_re <= _T_2618_re;
    _T_2619_im <= _T_2618_im;
    _T_2620_re <= _T_2619_re;
    _T_2620_im <= _T_2619_im;
    _T_2621_re <= _T_2620_re;
    _T_2621_im <= _T_2620_im;
    _T_2622_re <= _T_2621_re;
    _T_2622_im <= _T_2621_im;
    _T_2623_re <= _T_2622_re;
    _T_2623_im <= _T_2622_im;
    _T_2624_re <= _T_2623_re;
    _T_2624_im <= _T_2623_im;
    _T_2625_re <= _T_2624_re;
    _T_2625_im <= _T_2624_im;
    _T_2626_re <= _T_2625_re;
    _T_2626_im <= _T_2625_im;
    _T_2627_re <= _T_2626_re;
    _T_2627_im <= _T_2626_im;
    _T_2628_re <= _T_2627_re;
    _T_2628_im <= _T_2627_im;
    _T_2629_re <= _T_2628_re;
    _T_2629_im <= _T_2628_im;
    _T_2630_re <= _T_2629_re;
    _T_2630_im <= _T_2629_im;
    _T_2631_re <= _T_2630_re;
    _T_2631_im <= _T_2630_im;
    _T_2632_re <= _T_2631_re;
    _T_2632_im <= _T_2631_im;
    _T_2633_re <= _T_2632_re;
    _T_2633_im <= _T_2632_im;
    _T_2634_re <= _T_2633_re;
    _T_2634_im <= _T_2633_im;
    _T_2635_re <= _T_2634_re;
    _T_2635_im <= _T_2634_im;
    _T_2636_re <= _T_2635_re;
    _T_2636_im <= _T_2635_im;
    _T_2637_re <= _T_2636_re;
    _T_2637_im <= _T_2636_im;
    _T_2638_re <= _T_2637_re;
    _T_2638_im <= _T_2637_im;
    _T_2639_re <= _T_2638_re;
    _T_2639_im <= _T_2638_im;
    _T_2640_re <= _T_2639_re;
    _T_2640_im <= _T_2639_im;
    _T_2641_re <= _T_2640_re;
    _T_2641_im <= _T_2640_im;
    _T_2642_re <= _T_2641_re;
    _T_2642_im <= _T_2641_im;
    _T_2643_re <= _T_2642_re;
    _T_2643_im <= _T_2642_im;
    _T_2644_re <= _T_2643_re;
    _T_2644_im <= _T_2643_im;
    _T_2645_re <= _T_2644_re;
    _T_2645_im <= _T_2644_im;
    _T_2646_re <= _T_2645_re;
    _T_2646_im <= _T_2645_im;
    _T_2647_re <= _T_2646_re;
    _T_2647_im <= _T_2646_im;
    _T_2648_re <= _T_2647_re;
    _T_2648_im <= _T_2647_im;
    _T_2649_re <= _T_2648_re;
    _T_2649_im <= _T_2648_im;
    _T_2650_re <= _T_2649_re;
    _T_2650_im <= _T_2649_im;
    _T_2651_re <= _T_2650_re;
    _T_2651_im <= _T_2650_im;
    _T_2652_re <= _T_2651_re;
    _T_2652_im <= _T_2651_im;
    _T_2653_re <= _T_2652_re;
    _T_2653_im <= _T_2652_im;
    _T_2654_re <= _T_2653_re;
    _T_2654_im <= _T_2653_im;
    _T_2655_re <= _T_2654_re;
    _T_2655_im <= _T_2654_im;
    _T_2656_re <= _T_2655_re;
    _T_2656_im <= _T_2655_im;
    _T_2657_re <= _T_2656_re;
    _T_2657_im <= _T_2656_im;
    _T_2658_re <= _T_2657_re;
    _T_2658_im <= _T_2657_im;
    _T_2659_re <= _T_2658_re;
    _T_2659_im <= _T_2658_im;
    _T_2660_re <= _T_2659_re;
    _T_2660_im <= _T_2659_im;
    _T_2661_re <= _T_2660_re;
    _T_2661_im <= _T_2660_im;
    _T_2662_re <= _T_2661_re;
    _T_2662_im <= _T_2661_im;
    _T_2663_re <= _T_2662_re;
    _T_2663_im <= _T_2662_im;
    _T_2664_re <= _T_2663_re;
    _T_2664_im <= _T_2663_im;
    _T_2665_re <= _T_2664_re;
    _T_2665_im <= _T_2664_im;
    _T_2666_re <= _T_2665_re;
    _T_2666_im <= _T_2665_im;
    _T_2667_re <= _T_2666_re;
    _T_2667_im <= _T_2666_im;
    _T_2668_re <= _T_2667_re;
    _T_2668_im <= _T_2667_im;
    _T_2669_re <= _T_2668_re;
    _T_2669_im <= _T_2668_im;
    _T_2670_re <= _T_2669_re;
    _T_2670_im <= _T_2669_im;
    _T_2671_re <= _T_2670_re;
    _T_2671_im <= _T_2670_im;
    _T_2672_re <= _T_2671_re;
    _T_2672_im <= _T_2671_im;
    _T_2673_re <= _T_2672_re;
    _T_2673_im <= _T_2672_im;
    _T_2674_re <= _T_2673_re;
    _T_2674_im <= _T_2673_im;
    _T_2675_re <= _T_2674_re;
    _T_2675_im <= _T_2674_im;
    _T_2676_re <= _T_2675_re;
    _T_2676_im <= _T_2675_im;
    _T_2677_re <= _T_2676_re;
    _T_2677_im <= _T_2676_im;
    _T_2678_re <= _T_2677_re;
    _T_2678_im <= _T_2677_im;
    _T_2679_re <= _T_2678_re;
    _T_2679_im <= _T_2678_im;
    _T_2680_re <= _T_2679_re;
    _T_2680_im <= _T_2679_im;
    _T_2681_re <= _T_2680_re;
    _T_2681_im <= _T_2680_im;
    _T_2682_re <= _T_2681_re;
    _T_2682_im <= _T_2681_im;
    _T_2683_re <= _T_2682_re;
    _T_2683_im <= _T_2682_im;
    _T_2684_re <= _T_2683_re;
    _T_2684_im <= _T_2683_im;
    _T_2685_re <= _T_2684_re;
    _T_2685_im <= _T_2684_im;
    _T_2686_re <= _T_2685_re;
    _T_2686_im <= _T_2685_im;
    _T_2687_re <= _T_2686_re;
    _T_2687_im <= _T_2686_im;
    _T_2688_re <= _T_2687_re;
    _T_2688_im <= _T_2687_im;
    _T_2689_re <= _T_2688_re;
    _T_2689_im <= _T_2688_im;
    _T_2690_re <= _T_2689_re;
    _T_2690_im <= _T_2689_im;
    _T_2691_re <= _T_2690_re;
    _T_2691_im <= _T_2690_im;
    _T_2692_re <= _T_2691_re;
    _T_2692_im <= _T_2691_im;
    _T_2693_re <= _T_2692_re;
    _T_2693_im <= _T_2692_im;
    _T_2694_re <= _T_2693_re;
    _T_2694_im <= _T_2693_im;
    _T_2695_re <= _T_2694_re;
    _T_2695_im <= _T_2694_im;
    _T_2696_re <= _T_2695_re;
    _T_2696_im <= _T_2695_im;
    _T_2697_re <= _T_2696_re;
    _T_2697_im <= _T_2696_im;
    _T_2698_re <= _T_2697_re;
    _T_2698_im <= _T_2697_im;
    _T_2699_re <= _T_2698_re;
    _T_2699_im <= _T_2698_im;
    _T_2700_re <= _T_2699_re;
    _T_2700_im <= _T_2699_im;
    _T_2701_re <= _T_2700_re;
    _T_2701_im <= _T_2700_im;
    _T_2702_re <= _T_2701_re;
    _T_2702_im <= _T_2701_im;
    _T_2703_re <= _T_2702_re;
    _T_2703_im <= _T_2702_im;
    _T_2704_re <= _T_2703_re;
    _T_2704_im <= _T_2703_im;
    _T_2705_re <= _T_2704_re;
    _T_2705_im <= _T_2704_im;
    _T_2706_re <= _T_2705_re;
    _T_2706_im <= _T_2705_im;
    _T_2707_re <= _T_2706_re;
    _T_2707_im <= _T_2706_im;
    _T_2708_re <= _T_2707_re;
    _T_2708_im <= _T_2707_im;
    _T_2709_re <= _T_2708_re;
    _T_2709_im <= _T_2708_im;
    _T_2710_re <= _T_2709_re;
    _T_2710_im <= _T_2709_im;
    _T_2711_re <= _T_2710_re;
    _T_2711_im <= _T_2710_im;
    _T_2712_re <= _T_2711_re;
    _T_2712_im <= _T_2711_im;
    _T_2713_re <= _T_2712_re;
    _T_2713_im <= _T_2712_im;
    _T_2714_re <= _T_2713_re;
    _T_2714_im <= _T_2713_im;
    _T_2715_re <= _T_2714_re;
    _T_2715_im <= _T_2714_im;
    _T_2716_re <= _T_2715_re;
    _T_2716_im <= _T_2715_im;
    _T_2717_re <= _T_2716_re;
    _T_2717_im <= _T_2716_im;
    _T_2718_re <= _T_2717_re;
    _T_2718_im <= _T_2717_im;
    _T_2719_re <= _T_2718_re;
    _T_2719_im <= _T_2718_im;
    _T_2720_re <= _T_2719_re;
    _T_2720_im <= _T_2719_im;
    _T_2721_re <= _T_2720_re;
    _T_2721_im <= _T_2720_im;
    _T_2722_re <= _T_2721_re;
    _T_2722_im <= _T_2721_im;
    _T_2723_re <= _T_2722_re;
    _T_2723_im <= _T_2722_im;
    _T_2724_re <= _T_2723_re;
    _T_2724_im <= _T_2723_im;
    _T_2725_re <= _T_2724_re;
    _T_2725_im <= _T_2724_im;
    _T_2726_re <= _T_2725_re;
    _T_2726_im <= _T_2725_im;
    _T_2727_re <= _T_2726_re;
    _T_2727_im <= _T_2726_im;
    _T_2728_re <= _T_2727_re;
    _T_2728_im <= _T_2727_im;
    _T_2729_re <= _T_2728_re;
    _T_2729_im <= _T_2728_im;
    _T_2730_re <= _T_2729_re;
    _T_2730_im <= _T_2729_im;
    _T_2731_re <= _T_2730_re;
    _T_2731_im <= _T_2730_im;
    _T_2732_re <= _T_2731_re;
    _T_2732_im <= _T_2731_im;
    _T_2733_re <= _T_2732_re;
    _T_2733_im <= _T_2732_im;
    _T_2734_re <= _T_2733_re;
    _T_2734_im <= _T_2733_im;
    _T_2735_re <= _T_2734_re;
    _T_2735_im <= _T_2734_im;
    _T_2736_re <= _T_2735_re;
    _T_2736_im <= _T_2735_im;
    _T_2737_re <= _T_2736_re;
    _T_2737_im <= _T_2736_im;
    _T_2738_re <= _T_2737_re;
    _T_2738_im <= _T_2737_im;
    _T_2739_re <= _T_2738_re;
    _T_2739_im <= _T_2738_im;
    _T_2740_re <= _T_2739_re;
    _T_2740_im <= _T_2739_im;
    _T_2741_re <= _T_2740_re;
    _T_2741_im <= _T_2740_im;
    _T_2742_re <= _T_2741_re;
    _T_2742_im <= _T_2741_im;
    _T_2743_re <= _T_2742_re;
    _T_2743_im <= _T_2742_im;
    _T_2744_re <= _T_2743_re;
    _T_2744_im <= _T_2743_im;
    _T_2745_re <= _T_2744_re;
    _T_2745_im <= _T_2744_im;
    _T_2746_re <= _T_2745_re;
    _T_2746_im <= _T_2745_im;
    _T_2747_re <= _T_2746_re;
    _T_2747_im <= _T_2746_im;
    _T_2748_re <= _T_2747_re;
    _T_2748_im <= _T_2747_im;
    _T_2749_re <= _T_2748_re;
    _T_2749_im <= _T_2748_im;
    _T_2750_re <= _T_2749_re;
    _T_2750_im <= _T_2749_im;
    _T_2751_re <= _T_2750_re;
    _T_2751_im <= _T_2750_im;
    _T_2752_re <= _T_2751_re;
    _T_2752_im <= _T_2751_im;
    _T_2753_re <= _T_2752_re;
    _T_2753_im <= _T_2752_im;
    _T_2754_re <= _T_2753_re;
    _T_2754_im <= _T_2753_im;
    _T_2755_re <= _T_2754_re;
    _T_2755_im <= _T_2754_im;
    _T_2756_re <= _T_2755_re;
    _T_2756_im <= _T_2755_im;
    _T_2757_re <= _T_2756_re;
    _T_2757_im <= _T_2756_im;
    _T_2758_re <= _T_2757_re;
    _T_2758_im <= _T_2757_im;
    _T_2759_re <= _T_2758_re;
    _T_2759_im <= _T_2758_im;
    _T_2760_re <= _T_2759_re;
    _T_2760_im <= _T_2759_im;
    _T_2761_re <= _T_2760_re;
    _T_2761_im <= _T_2760_im;
    _T_2762_re <= _T_2761_re;
    _T_2762_im <= _T_2761_im;
    _T_2765_re <= Butterfly_2_io_out2_re;
    _T_2765_im <= Butterfly_2_io_out2_im;
    _T_2766_re <= _T_2765_re;
    _T_2766_im <= _T_2765_im;
    _T_2767_re <= _T_2766_re;
    _T_2767_im <= _T_2766_im;
    _T_2768_re <= _T_2767_re;
    _T_2768_im <= _T_2767_im;
    _T_2769_re <= _T_2768_re;
    _T_2769_im <= _T_2768_im;
    _T_2770_re <= _T_2769_re;
    _T_2770_im <= _T_2769_im;
    _T_2771_re <= _T_2770_re;
    _T_2771_im <= _T_2770_im;
    _T_2772_re <= _T_2771_re;
    _T_2772_im <= _T_2771_im;
    _T_2773_re <= _T_2772_re;
    _T_2773_im <= _T_2772_im;
    _T_2774_re <= _T_2773_re;
    _T_2774_im <= _T_2773_im;
    _T_2775_re <= _T_2774_re;
    _T_2775_im <= _T_2774_im;
    _T_2776_re <= _T_2775_re;
    _T_2776_im <= _T_2775_im;
    _T_2777_re <= _T_2776_re;
    _T_2777_im <= _T_2776_im;
    _T_2778_re <= _T_2777_re;
    _T_2778_im <= _T_2777_im;
    _T_2779_re <= _T_2778_re;
    _T_2779_im <= _T_2778_im;
    _T_2780_re <= _T_2779_re;
    _T_2780_im <= _T_2779_im;
    _T_2781_re <= _T_2780_re;
    _T_2781_im <= _T_2780_im;
    _T_2782_re <= _T_2781_re;
    _T_2782_im <= _T_2781_im;
    _T_2783_re <= _T_2782_re;
    _T_2783_im <= _T_2782_im;
    _T_2784_re <= _T_2783_re;
    _T_2784_im <= _T_2783_im;
    _T_2785_re <= _T_2784_re;
    _T_2785_im <= _T_2784_im;
    _T_2786_re <= _T_2785_re;
    _T_2786_im <= _T_2785_im;
    _T_2787_re <= _T_2786_re;
    _T_2787_im <= _T_2786_im;
    _T_2788_re <= _T_2787_re;
    _T_2788_im <= _T_2787_im;
    _T_2789_re <= _T_2788_re;
    _T_2789_im <= _T_2788_im;
    _T_2790_re <= _T_2789_re;
    _T_2790_im <= _T_2789_im;
    _T_2791_re <= _T_2790_re;
    _T_2791_im <= _T_2790_im;
    _T_2792_re <= _T_2791_re;
    _T_2792_im <= _T_2791_im;
    _T_2793_re <= _T_2792_re;
    _T_2793_im <= _T_2792_im;
    _T_2794_re <= _T_2793_re;
    _T_2794_im <= _T_2793_im;
    _T_2795_re <= _T_2794_re;
    _T_2795_im <= _T_2794_im;
    _T_2796_re <= _T_2795_re;
    _T_2796_im <= _T_2795_im;
    _T_2797_re <= _T_2796_re;
    _T_2797_im <= _T_2796_im;
    _T_2798_re <= _T_2797_re;
    _T_2798_im <= _T_2797_im;
    _T_2799_re <= _T_2798_re;
    _T_2799_im <= _T_2798_im;
    _T_2800_re <= _T_2799_re;
    _T_2800_im <= _T_2799_im;
    _T_2801_re <= _T_2800_re;
    _T_2801_im <= _T_2800_im;
    _T_2802_re <= _T_2801_re;
    _T_2802_im <= _T_2801_im;
    _T_2803_re <= _T_2802_re;
    _T_2803_im <= _T_2802_im;
    _T_2804_re <= _T_2803_re;
    _T_2804_im <= _T_2803_im;
    _T_2805_re <= _T_2804_re;
    _T_2805_im <= _T_2804_im;
    _T_2806_re <= _T_2805_re;
    _T_2806_im <= _T_2805_im;
    _T_2807_re <= _T_2806_re;
    _T_2807_im <= _T_2806_im;
    _T_2808_re <= _T_2807_re;
    _T_2808_im <= _T_2807_im;
    _T_2809_re <= _T_2808_re;
    _T_2809_im <= _T_2808_im;
    _T_2810_re <= _T_2809_re;
    _T_2810_im <= _T_2809_im;
    _T_2811_re <= _T_2810_re;
    _T_2811_im <= _T_2810_im;
    _T_2812_re <= _T_2811_re;
    _T_2812_im <= _T_2811_im;
    _T_2813_re <= _T_2812_re;
    _T_2813_im <= _T_2812_im;
    _T_2814_re <= _T_2813_re;
    _T_2814_im <= _T_2813_im;
    _T_2815_re <= _T_2814_re;
    _T_2815_im <= _T_2814_im;
    _T_2816_re <= _T_2815_re;
    _T_2816_im <= _T_2815_im;
    _T_2817_re <= _T_2816_re;
    _T_2817_im <= _T_2816_im;
    _T_2818_re <= _T_2817_re;
    _T_2818_im <= _T_2817_im;
    _T_2819_re <= _T_2818_re;
    _T_2819_im <= _T_2818_im;
    _T_2820_re <= _T_2819_re;
    _T_2820_im <= _T_2819_im;
    _T_2821_re <= _T_2820_re;
    _T_2821_im <= _T_2820_im;
    _T_2822_re <= _T_2821_re;
    _T_2822_im <= _T_2821_im;
    _T_2823_re <= _T_2822_re;
    _T_2823_im <= _T_2822_im;
    _T_2824_re <= _T_2823_re;
    _T_2824_im <= _T_2823_im;
    _T_2825_re <= _T_2824_re;
    _T_2825_im <= _T_2824_im;
    _T_2826_re <= _T_2825_re;
    _T_2826_im <= _T_2825_im;
    _T_2827_re <= _T_2826_re;
    _T_2827_im <= _T_2826_im;
    _T_2828_re <= _T_2827_re;
    _T_2828_im <= _T_2827_im;
    _T_2829_re <= _T_2828_re;
    _T_2829_im <= _T_2828_im;
    _T_2830_re <= _T_2829_re;
    _T_2830_im <= _T_2829_im;
    _T_2831_re <= _T_2830_re;
    _T_2831_im <= _T_2830_im;
    _T_2832_re <= _T_2831_re;
    _T_2832_im <= _T_2831_im;
    _T_2833_re <= _T_2832_re;
    _T_2833_im <= _T_2832_im;
    _T_2834_re <= _T_2833_re;
    _T_2834_im <= _T_2833_im;
    _T_2835_re <= _T_2834_re;
    _T_2835_im <= _T_2834_im;
    _T_2836_re <= _T_2835_re;
    _T_2836_im <= _T_2835_im;
    _T_2837_re <= _T_2836_re;
    _T_2837_im <= _T_2836_im;
    _T_2838_re <= _T_2837_re;
    _T_2838_im <= _T_2837_im;
    _T_2839_re <= _T_2838_re;
    _T_2839_im <= _T_2838_im;
    _T_2840_re <= _T_2839_re;
    _T_2840_im <= _T_2839_im;
    _T_2841_re <= _T_2840_re;
    _T_2841_im <= _T_2840_im;
    _T_2842_re <= _T_2841_re;
    _T_2842_im <= _T_2841_im;
    _T_2843_re <= _T_2842_re;
    _T_2843_im <= _T_2842_im;
    _T_2844_re <= _T_2843_re;
    _T_2844_im <= _T_2843_im;
    _T_2845_re <= _T_2844_re;
    _T_2845_im <= _T_2844_im;
    _T_2846_re <= _T_2845_re;
    _T_2846_im <= _T_2845_im;
    _T_2847_re <= _T_2846_re;
    _T_2847_im <= _T_2846_im;
    _T_2848_re <= _T_2847_re;
    _T_2848_im <= _T_2847_im;
    _T_2849_re <= _T_2848_re;
    _T_2849_im <= _T_2848_im;
    _T_2850_re <= _T_2849_re;
    _T_2850_im <= _T_2849_im;
    _T_2851_re <= _T_2850_re;
    _T_2851_im <= _T_2850_im;
    _T_2852_re <= _T_2851_re;
    _T_2852_im <= _T_2851_im;
    _T_2853_re <= _T_2852_re;
    _T_2853_im <= _T_2852_im;
    _T_2854_re <= _T_2853_re;
    _T_2854_im <= _T_2853_im;
    _T_2855_re <= _T_2854_re;
    _T_2855_im <= _T_2854_im;
    _T_2856_re <= _T_2855_re;
    _T_2856_im <= _T_2855_im;
    _T_2857_re <= _T_2856_re;
    _T_2857_im <= _T_2856_im;
    _T_2858_re <= _T_2857_re;
    _T_2858_im <= _T_2857_im;
    _T_2859_re <= _T_2858_re;
    _T_2859_im <= _T_2858_im;
    _T_2860_re <= _T_2859_re;
    _T_2860_im <= _T_2859_im;
    _T_2861_re <= _T_2860_re;
    _T_2861_im <= _T_2860_im;
    _T_2862_re <= _T_2861_re;
    _T_2862_im <= _T_2861_im;
    _T_2863_re <= _T_2862_re;
    _T_2863_im <= _T_2862_im;
    _T_2864_re <= _T_2863_re;
    _T_2864_im <= _T_2863_im;
    _T_2865_re <= _T_2864_re;
    _T_2865_im <= _T_2864_im;
    _T_2866_re <= _T_2865_re;
    _T_2866_im <= _T_2865_im;
    _T_2867_re <= _T_2866_re;
    _T_2867_im <= _T_2866_im;
    _T_2868_re <= _T_2867_re;
    _T_2868_im <= _T_2867_im;
    _T_2869_re <= _T_2868_re;
    _T_2869_im <= _T_2868_im;
    _T_2870_re <= _T_2869_re;
    _T_2870_im <= _T_2869_im;
    _T_2871_re <= _T_2870_re;
    _T_2871_im <= _T_2870_im;
    _T_2872_re <= _T_2871_re;
    _T_2872_im <= _T_2871_im;
    _T_2873_re <= _T_2872_re;
    _T_2873_im <= _T_2872_im;
    _T_2874_re <= _T_2873_re;
    _T_2874_im <= _T_2873_im;
    _T_2875_re <= _T_2874_re;
    _T_2875_im <= _T_2874_im;
    _T_2876_re <= _T_2875_re;
    _T_2876_im <= _T_2875_im;
    _T_2877_re <= _T_2876_re;
    _T_2877_im <= _T_2876_im;
    _T_2878_re <= _T_2877_re;
    _T_2878_im <= _T_2877_im;
    _T_2879_re <= _T_2878_re;
    _T_2879_im <= _T_2878_im;
    _T_2880_re <= _T_2879_re;
    _T_2880_im <= _T_2879_im;
    _T_2881_re <= _T_2880_re;
    _T_2881_im <= _T_2880_im;
    _T_2882_re <= _T_2881_re;
    _T_2882_im <= _T_2881_im;
    _T_2883_re <= _T_2882_re;
    _T_2883_im <= _T_2882_im;
    _T_2884_re <= _T_2883_re;
    _T_2884_im <= _T_2883_im;
    _T_2885_re <= _T_2884_re;
    _T_2885_im <= _T_2884_im;
    _T_2886_re <= _T_2885_re;
    _T_2886_im <= _T_2885_im;
    _T_2887_re <= _T_2886_re;
    _T_2887_im <= _T_2886_im;
    _T_2888_re <= _T_2887_re;
    _T_2888_im <= _T_2887_im;
    _T_2889_re <= _T_2888_re;
    _T_2889_im <= _T_2888_im;
    _T_2890_re <= _T_2889_re;
    _T_2890_im <= _T_2889_im;
    _T_2891_re <= _T_2890_re;
    _T_2891_im <= _T_2890_im;
    _T_2892_re <= _T_2891_re;
    _T_2892_im <= _T_2891_im;
    _T_2902_re <= Switch_2_io_out1_re;
    _T_2902_im <= Switch_2_io_out1_im;
    _T_2903_re <= _T_2902_re;
    _T_2903_im <= _T_2902_im;
    _T_2904_re <= _T_2903_re;
    _T_2904_im <= _T_2903_im;
    _T_2905_re <= _T_2904_re;
    _T_2905_im <= _T_2904_im;
    _T_2906_re <= _T_2905_re;
    _T_2906_im <= _T_2905_im;
    _T_2907_re <= _T_2906_re;
    _T_2907_im <= _T_2906_im;
    _T_2908_re <= _T_2907_re;
    _T_2908_im <= _T_2907_im;
    _T_2909_re <= _T_2908_re;
    _T_2909_im <= _T_2908_im;
    _T_2910_re <= _T_2909_re;
    _T_2910_im <= _T_2909_im;
    _T_2911_re <= _T_2910_re;
    _T_2911_im <= _T_2910_im;
    _T_2912_re <= _T_2911_re;
    _T_2912_im <= _T_2911_im;
    _T_2913_re <= _T_2912_re;
    _T_2913_im <= _T_2912_im;
    _T_2914_re <= _T_2913_re;
    _T_2914_im <= _T_2913_im;
    _T_2915_re <= _T_2914_re;
    _T_2915_im <= _T_2914_im;
    _T_2916_re <= _T_2915_re;
    _T_2916_im <= _T_2915_im;
    _T_2917_re <= _T_2916_re;
    _T_2917_im <= _T_2916_im;
    _T_2918_re <= _T_2917_re;
    _T_2918_im <= _T_2917_im;
    _T_2919_re <= _T_2918_re;
    _T_2919_im <= _T_2918_im;
    _T_2920_re <= _T_2919_re;
    _T_2920_im <= _T_2919_im;
    _T_2921_re <= _T_2920_re;
    _T_2921_im <= _T_2920_im;
    _T_2922_re <= _T_2921_re;
    _T_2922_im <= _T_2921_im;
    _T_2923_re <= _T_2922_re;
    _T_2923_im <= _T_2922_im;
    _T_2924_re <= _T_2923_re;
    _T_2924_im <= _T_2923_im;
    _T_2925_re <= _T_2924_re;
    _T_2925_im <= _T_2924_im;
    _T_2926_re <= _T_2925_re;
    _T_2926_im <= _T_2925_im;
    _T_2927_re <= _T_2926_re;
    _T_2927_im <= _T_2926_im;
    _T_2928_re <= _T_2927_re;
    _T_2928_im <= _T_2927_im;
    _T_2929_re <= _T_2928_re;
    _T_2929_im <= _T_2928_im;
    _T_2930_re <= _T_2929_re;
    _T_2930_im <= _T_2929_im;
    _T_2931_re <= _T_2930_re;
    _T_2931_im <= _T_2930_im;
    _T_2932_re <= _T_2931_re;
    _T_2932_im <= _T_2931_im;
    _T_2933_re <= _T_2932_re;
    _T_2933_im <= _T_2932_im;
    _T_2934_re <= _T_2933_re;
    _T_2934_im <= _T_2933_im;
    _T_2935_re <= _T_2934_re;
    _T_2935_im <= _T_2934_im;
    _T_2936_re <= _T_2935_re;
    _T_2936_im <= _T_2935_im;
    _T_2937_re <= _T_2936_re;
    _T_2937_im <= _T_2936_im;
    _T_2938_re <= _T_2937_re;
    _T_2938_im <= _T_2937_im;
    _T_2939_re <= _T_2938_re;
    _T_2939_im <= _T_2938_im;
    _T_2940_re <= _T_2939_re;
    _T_2940_im <= _T_2939_im;
    _T_2941_re <= _T_2940_re;
    _T_2941_im <= _T_2940_im;
    _T_2942_re <= _T_2941_re;
    _T_2942_im <= _T_2941_im;
    _T_2943_re <= _T_2942_re;
    _T_2943_im <= _T_2942_im;
    _T_2944_re <= _T_2943_re;
    _T_2944_im <= _T_2943_im;
    _T_2945_re <= _T_2944_re;
    _T_2945_im <= _T_2944_im;
    _T_2946_re <= _T_2945_re;
    _T_2946_im <= _T_2945_im;
    _T_2947_re <= _T_2946_re;
    _T_2947_im <= _T_2946_im;
    _T_2948_re <= _T_2947_re;
    _T_2948_im <= _T_2947_im;
    _T_2949_re <= _T_2948_re;
    _T_2949_im <= _T_2948_im;
    _T_2950_re <= _T_2949_re;
    _T_2950_im <= _T_2949_im;
    _T_2951_re <= _T_2950_re;
    _T_2951_im <= _T_2950_im;
    _T_2952_re <= _T_2951_re;
    _T_2952_im <= _T_2951_im;
    _T_2953_re <= _T_2952_re;
    _T_2953_im <= _T_2952_im;
    _T_2954_re <= _T_2953_re;
    _T_2954_im <= _T_2953_im;
    _T_2955_re <= _T_2954_re;
    _T_2955_im <= _T_2954_im;
    _T_2956_re <= _T_2955_re;
    _T_2956_im <= _T_2955_im;
    _T_2957_re <= _T_2956_re;
    _T_2957_im <= _T_2956_im;
    _T_2958_re <= _T_2957_re;
    _T_2958_im <= _T_2957_im;
    _T_2959_re <= _T_2958_re;
    _T_2959_im <= _T_2958_im;
    _T_2960_re <= _T_2959_re;
    _T_2960_im <= _T_2959_im;
    _T_2961_re <= _T_2960_re;
    _T_2961_im <= _T_2960_im;
    _T_2962_re <= _T_2961_re;
    _T_2962_im <= _T_2961_im;
    _T_2963_re <= _T_2962_re;
    _T_2963_im <= _T_2962_im;
    _T_2964_re <= _T_2963_re;
    _T_2964_im <= _T_2963_im;
    _T_2965_re <= _T_2964_re;
    _T_2965_im <= _T_2964_im;
    _T_2966_re <= _T_2965_re;
    _T_2966_im <= _T_2965_im;
    _T_2967_re <= _T_2966_re;
    _T_2967_im <= _T_2966_im;
    _T_2968_re <= _T_2967_re;
    _T_2968_im <= _T_2967_im;
    _T_2969_re <= _T_2968_re;
    _T_2969_im <= _T_2968_im;
    _T_2970_re <= _T_2969_re;
    _T_2970_im <= _T_2969_im;
    _T_2971_re <= _T_2970_re;
    _T_2971_im <= _T_2970_im;
    _T_2972_re <= _T_2971_re;
    _T_2972_im <= _T_2971_im;
    _T_2973_re <= _T_2972_re;
    _T_2973_im <= _T_2972_im;
    _T_2974_re <= _T_2973_re;
    _T_2974_im <= _T_2973_im;
    _T_2975_re <= _T_2974_re;
    _T_2975_im <= _T_2974_im;
    _T_2976_re <= _T_2975_re;
    _T_2976_im <= _T_2975_im;
    _T_2977_re <= _T_2976_re;
    _T_2977_im <= _T_2976_im;
    _T_2978_re <= _T_2977_re;
    _T_2978_im <= _T_2977_im;
    _T_2979_re <= _T_2978_re;
    _T_2979_im <= _T_2978_im;
    _T_2980_re <= _T_2979_re;
    _T_2980_im <= _T_2979_im;
    _T_2981_re <= _T_2980_re;
    _T_2981_im <= _T_2980_im;
    _T_2982_re <= _T_2981_re;
    _T_2982_im <= _T_2981_im;
    _T_2983_re <= _T_2982_re;
    _T_2983_im <= _T_2982_im;
    _T_2984_re <= _T_2983_re;
    _T_2984_im <= _T_2983_im;
    _T_2985_re <= _T_2984_re;
    _T_2985_im <= _T_2984_im;
    _T_2986_re <= _T_2985_re;
    _T_2986_im <= _T_2985_im;
    _T_2987_re <= _T_2986_re;
    _T_2987_im <= _T_2986_im;
    _T_2988_re <= _T_2987_re;
    _T_2988_im <= _T_2987_im;
    _T_2989_re <= _T_2988_re;
    _T_2989_im <= _T_2988_im;
    _T_2990_re <= _T_2989_re;
    _T_2990_im <= _T_2989_im;
    _T_2991_re <= _T_2990_re;
    _T_2991_im <= _T_2990_im;
    _T_2992_re <= _T_2991_re;
    _T_2992_im <= _T_2991_im;
    _T_2993_re <= _T_2992_re;
    _T_2993_im <= _T_2992_im;
    _T_2994_re <= _T_2993_re;
    _T_2994_im <= _T_2993_im;
    _T_2995_re <= _T_2994_re;
    _T_2995_im <= _T_2994_im;
    _T_2996_re <= _T_2995_re;
    _T_2996_im <= _T_2995_im;
    _T_2997_re <= _T_2996_re;
    _T_2997_im <= _T_2996_im;
    _T_2998_re <= _T_2997_re;
    _T_2998_im <= _T_2997_im;
    _T_2999_re <= _T_2998_re;
    _T_2999_im <= _T_2998_im;
    _T_3000_re <= _T_2999_re;
    _T_3000_im <= _T_2999_im;
    _T_3001_re <= _T_3000_re;
    _T_3001_im <= _T_3000_im;
    _T_3002_re <= _T_3001_re;
    _T_3002_im <= _T_3001_im;
    _T_3003_re <= _T_3002_re;
    _T_3003_im <= _T_3002_im;
    _T_3004_re <= _T_3003_re;
    _T_3004_im <= _T_3003_im;
    _T_3005_re <= _T_3004_re;
    _T_3005_im <= _T_3004_im;
    _T_3006_re <= _T_3005_re;
    _T_3006_im <= _T_3005_im;
    _T_3007_re <= _T_3006_re;
    _T_3007_im <= _T_3006_im;
    _T_3008_re <= _T_3007_re;
    _T_3008_im <= _T_3007_im;
    _T_3009_re <= _T_3008_re;
    _T_3009_im <= _T_3008_im;
    _T_3010_re <= _T_3009_re;
    _T_3010_im <= _T_3009_im;
    _T_3011_re <= _T_3010_re;
    _T_3011_im <= _T_3010_im;
    _T_3012_re <= _T_3011_re;
    _T_3012_im <= _T_3011_im;
    _T_3013_re <= _T_3012_re;
    _T_3013_im <= _T_3012_im;
    _T_3014_re <= _T_3013_re;
    _T_3014_im <= _T_3013_im;
    _T_3015_re <= _T_3014_re;
    _T_3015_im <= _T_3014_im;
    _T_3016_re <= _T_3015_re;
    _T_3016_im <= _T_3015_im;
    _T_3017_re <= _T_3016_re;
    _T_3017_im <= _T_3016_im;
    _T_3018_re <= _T_3017_re;
    _T_3018_im <= _T_3017_im;
    _T_3019_re <= _T_3018_re;
    _T_3019_im <= _T_3018_im;
    _T_3020_re <= _T_3019_re;
    _T_3020_im <= _T_3019_im;
    _T_3021_re <= _T_3020_re;
    _T_3021_im <= _T_3020_im;
    _T_3022_re <= _T_3021_re;
    _T_3022_im <= _T_3021_im;
    _T_3023_re <= _T_3022_re;
    _T_3023_im <= _T_3022_im;
    _T_3024_re <= _T_3023_re;
    _T_3024_im <= _T_3023_im;
    _T_3025_re <= _T_3024_re;
    _T_3025_im <= _T_3024_im;
    _T_3026_re <= _T_3025_re;
    _T_3026_im <= _T_3025_im;
    _T_3027_re <= _T_3026_re;
    _T_3027_im <= _T_3026_im;
    _T_3028_re <= _T_3027_re;
    _T_3028_im <= _T_3027_im;
    _T_3029_re <= _T_3028_re;
    _T_3029_im <= _T_3028_im;
    _T_3032_re <= Butterfly_3_io_out2_re;
    _T_3032_im <= Butterfly_3_io_out2_im;
    _T_3033_re <= _T_3032_re;
    _T_3033_im <= _T_3032_im;
    _T_3034_re <= _T_3033_re;
    _T_3034_im <= _T_3033_im;
    _T_3035_re <= _T_3034_re;
    _T_3035_im <= _T_3034_im;
    _T_3036_re <= _T_3035_re;
    _T_3036_im <= _T_3035_im;
    _T_3037_re <= _T_3036_re;
    _T_3037_im <= _T_3036_im;
    _T_3038_re <= _T_3037_re;
    _T_3038_im <= _T_3037_im;
    _T_3039_re <= _T_3038_re;
    _T_3039_im <= _T_3038_im;
    _T_3040_re <= _T_3039_re;
    _T_3040_im <= _T_3039_im;
    _T_3041_re <= _T_3040_re;
    _T_3041_im <= _T_3040_im;
    _T_3042_re <= _T_3041_re;
    _T_3042_im <= _T_3041_im;
    _T_3043_re <= _T_3042_re;
    _T_3043_im <= _T_3042_im;
    _T_3044_re <= _T_3043_re;
    _T_3044_im <= _T_3043_im;
    _T_3045_re <= _T_3044_re;
    _T_3045_im <= _T_3044_im;
    _T_3046_re <= _T_3045_re;
    _T_3046_im <= _T_3045_im;
    _T_3047_re <= _T_3046_re;
    _T_3047_im <= _T_3046_im;
    _T_3048_re <= _T_3047_re;
    _T_3048_im <= _T_3047_im;
    _T_3049_re <= _T_3048_re;
    _T_3049_im <= _T_3048_im;
    _T_3050_re <= _T_3049_re;
    _T_3050_im <= _T_3049_im;
    _T_3051_re <= _T_3050_re;
    _T_3051_im <= _T_3050_im;
    _T_3052_re <= _T_3051_re;
    _T_3052_im <= _T_3051_im;
    _T_3053_re <= _T_3052_re;
    _T_3053_im <= _T_3052_im;
    _T_3054_re <= _T_3053_re;
    _T_3054_im <= _T_3053_im;
    _T_3055_re <= _T_3054_re;
    _T_3055_im <= _T_3054_im;
    _T_3056_re <= _T_3055_re;
    _T_3056_im <= _T_3055_im;
    _T_3057_re <= _T_3056_re;
    _T_3057_im <= _T_3056_im;
    _T_3058_re <= _T_3057_re;
    _T_3058_im <= _T_3057_im;
    _T_3059_re <= _T_3058_re;
    _T_3059_im <= _T_3058_im;
    _T_3060_re <= _T_3059_re;
    _T_3060_im <= _T_3059_im;
    _T_3061_re <= _T_3060_re;
    _T_3061_im <= _T_3060_im;
    _T_3062_re <= _T_3061_re;
    _T_3062_im <= _T_3061_im;
    _T_3063_re <= _T_3062_re;
    _T_3063_im <= _T_3062_im;
    _T_3064_re <= _T_3063_re;
    _T_3064_im <= _T_3063_im;
    _T_3065_re <= _T_3064_re;
    _T_3065_im <= _T_3064_im;
    _T_3066_re <= _T_3065_re;
    _T_3066_im <= _T_3065_im;
    _T_3067_re <= _T_3066_re;
    _T_3067_im <= _T_3066_im;
    _T_3068_re <= _T_3067_re;
    _T_3068_im <= _T_3067_im;
    _T_3069_re <= _T_3068_re;
    _T_3069_im <= _T_3068_im;
    _T_3070_re <= _T_3069_re;
    _T_3070_im <= _T_3069_im;
    _T_3071_re <= _T_3070_re;
    _T_3071_im <= _T_3070_im;
    _T_3072_re <= _T_3071_re;
    _T_3072_im <= _T_3071_im;
    _T_3073_re <= _T_3072_re;
    _T_3073_im <= _T_3072_im;
    _T_3074_re <= _T_3073_re;
    _T_3074_im <= _T_3073_im;
    _T_3075_re <= _T_3074_re;
    _T_3075_im <= _T_3074_im;
    _T_3076_re <= _T_3075_re;
    _T_3076_im <= _T_3075_im;
    _T_3077_re <= _T_3076_re;
    _T_3077_im <= _T_3076_im;
    _T_3078_re <= _T_3077_re;
    _T_3078_im <= _T_3077_im;
    _T_3079_re <= _T_3078_re;
    _T_3079_im <= _T_3078_im;
    _T_3080_re <= _T_3079_re;
    _T_3080_im <= _T_3079_im;
    _T_3081_re <= _T_3080_re;
    _T_3081_im <= _T_3080_im;
    _T_3082_re <= _T_3081_re;
    _T_3082_im <= _T_3081_im;
    _T_3083_re <= _T_3082_re;
    _T_3083_im <= _T_3082_im;
    _T_3084_re <= _T_3083_re;
    _T_3084_im <= _T_3083_im;
    _T_3085_re <= _T_3084_re;
    _T_3085_im <= _T_3084_im;
    _T_3086_re <= _T_3085_re;
    _T_3086_im <= _T_3085_im;
    _T_3087_re <= _T_3086_re;
    _T_3087_im <= _T_3086_im;
    _T_3088_re <= _T_3087_re;
    _T_3088_im <= _T_3087_im;
    _T_3089_re <= _T_3088_re;
    _T_3089_im <= _T_3088_im;
    _T_3090_re <= _T_3089_re;
    _T_3090_im <= _T_3089_im;
    _T_3091_re <= _T_3090_re;
    _T_3091_im <= _T_3090_im;
    _T_3092_re <= _T_3091_re;
    _T_3092_im <= _T_3091_im;
    _T_3093_re <= _T_3092_re;
    _T_3093_im <= _T_3092_im;
    _T_3094_re <= _T_3093_re;
    _T_3094_im <= _T_3093_im;
    _T_3095_re <= _T_3094_re;
    _T_3095_im <= _T_3094_im;
    _T_3105_re <= Switch_3_io_out1_re;
    _T_3105_im <= Switch_3_io_out1_im;
    _T_3106_re <= _T_3105_re;
    _T_3106_im <= _T_3105_im;
    _T_3107_re <= _T_3106_re;
    _T_3107_im <= _T_3106_im;
    _T_3108_re <= _T_3107_re;
    _T_3108_im <= _T_3107_im;
    _T_3109_re <= _T_3108_re;
    _T_3109_im <= _T_3108_im;
    _T_3110_re <= _T_3109_re;
    _T_3110_im <= _T_3109_im;
    _T_3111_re <= _T_3110_re;
    _T_3111_im <= _T_3110_im;
    _T_3112_re <= _T_3111_re;
    _T_3112_im <= _T_3111_im;
    _T_3113_re <= _T_3112_re;
    _T_3113_im <= _T_3112_im;
    _T_3114_re <= _T_3113_re;
    _T_3114_im <= _T_3113_im;
    _T_3115_re <= _T_3114_re;
    _T_3115_im <= _T_3114_im;
    _T_3116_re <= _T_3115_re;
    _T_3116_im <= _T_3115_im;
    _T_3117_re <= _T_3116_re;
    _T_3117_im <= _T_3116_im;
    _T_3118_re <= _T_3117_re;
    _T_3118_im <= _T_3117_im;
    _T_3119_re <= _T_3118_re;
    _T_3119_im <= _T_3118_im;
    _T_3120_re <= _T_3119_re;
    _T_3120_im <= _T_3119_im;
    _T_3121_re <= _T_3120_re;
    _T_3121_im <= _T_3120_im;
    _T_3122_re <= _T_3121_re;
    _T_3122_im <= _T_3121_im;
    _T_3123_re <= _T_3122_re;
    _T_3123_im <= _T_3122_im;
    _T_3124_re <= _T_3123_re;
    _T_3124_im <= _T_3123_im;
    _T_3125_re <= _T_3124_re;
    _T_3125_im <= _T_3124_im;
    _T_3126_re <= _T_3125_re;
    _T_3126_im <= _T_3125_im;
    _T_3127_re <= _T_3126_re;
    _T_3127_im <= _T_3126_im;
    _T_3128_re <= _T_3127_re;
    _T_3128_im <= _T_3127_im;
    _T_3129_re <= _T_3128_re;
    _T_3129_im <= _T_3128_im;
    _T_3130_re <= _T_3129_re;
    _T_3130_im <= _T_3129_im;
    _T_3131_re <= _T_3130_re;
    _T_3131_im <= _T_3130_im;
    _T_3132_re <= _T_3131_re;
    _T_3132_im <= _T_3131_im;
    _T_3133_re <= _T_3132_re;
    _T_3133_im <= _T_3132_im;
    _T_3134_re <= _T_3133_re;
    _T_3134_im <= _T_3133_im;
    _T_3135_re <= _T_3134_re;
    _T_3135_im <= _T_3134_im;
    _T_3136_re <= _T_3135_re;
    _T_3136_im <= _T_3135_im;
    _T_3137_re <= _T_3136_re;
    _T_3137_im <= _T_3136_im;
    _T_3138_re <= _T_3137_re;
    _T_3138_im <= _T_3137_im;
    _T_3139_re <= _T_3138_re;
    _T_3139_im <= _T_3138_im;
    _T_3140_re <= _T_3139_re;
    _T_3140_im <= _T_3139_im;
    _T_3141_re <= _T_3140_re;
    _T_3141_im <= _T_3140_im;
    _T_3142_re <= _T_3141_re;
    _T_3142_im <= _T_3141_im;
    _T_3143_re <= _T_3142_re;
    _T_3143_im <= _T_3142_im;
    _T_3144_re <= _T_3143_re;
    _T_3144_im <= _T_3143_im;
    _T_3145_re <= _T_3144_re;
    _T_3145_im <= _T_3144_im;
    _T_3146_re <= _T_3145_re;
    _T_3146_im <= _T_3145_im;
    _T_3147_re <= _T_3146_re;
    _T_3147_im <= _T_3146_im;
    _T_3148_re <= _T_3147_re;
    _T_3148_im <= _T_3147_im;
    _T_3149_re <= _T_3148_re;
    _T_3149_im <= _T_3148_im;
    _T_3150_re <= _T_3149_re;
    _T_3150_im <= _T_3149_im;
    _T_3151_re <= _T_3150_re;
    _T_3151_im <= _T_3150_im;
    _T_3152_re <= _T_3151_re;
    _T_3152_im <= _T_3151_im;
    _T_3153_re <= _T_3152_re;
    _T_3153_im <= _T_3152_im;
    _T_3154_re <= _T_3153_re;
    _T_3154_im <= _T_3153_im;
    _T_3155_re <= _T_3154_re;
    _T_3155_im <= _T_3154_im;
    _T_3156_re <= _T_3155_re;
    _T_3156_im <= _T_3155_im;
    _T_3157_re <= _T_3156_re;
    _T_3157_im <= _T_3156_im;
    _T_3158_re <= _T_3157_re;
    _T_3158_im <= _T_3157_im;
    _T_3159_re <= _T_3158_re;
    _T_3159_im <= _T_3158_im;
    _T_3160_re <= _T_3159_re;
    _T_3160_im <= _T_3159_im;
    _T_3161_re <= _T_3160_re;
    _T_3161_im <= _T_3160_im;
    _T_3162_re <= _T_3161_re;
    _T_3162_im <= _T_3161_im;
    _T_3163_re <= _T_3162_re;
    _T_3163_im <= _T_3162_im;
    _T_3164_re <= _T_3163_re;
    _T_3164_im <= _T_3163_im;
    _T_3165_re <= _T_3164_re;
    _T_3165_im <= _T_3164_im;
    _T_3166_re <= _T_3165_re;
    _T_3166_im <= _T_3165_im;
    _T_3167_re <= _T_3166_re;
    _T_3167_im <= _T_3166_im;
    _T_3168_re <= _T_3167_re;
    _T_3168_im <= _T_3167_im;
    _T_3171_re <= Butterfly_4_io_out2_re;
    _T_3171_im <= Butterfly_4_io_out2_im;
    _T_3172_re <= _T_3171_re;
    _T_3172_im <= _T_3171_im;
    _T_3173_re <= _T_3172_re;
    _T_3173_im <= _T_3172_im;
    _T_3174_re <= _T_3173_re;
    _T_3174_im <= _T_3173_im;
    _T_3175_re <= _T_3174_re;
    _T_3175_im <= _T_3174_im;
    _T_3176_re <= _T_3175_re;
    _T_3176_im <= _T_3175_im;
    _T_3177_re <= _T_3176_re;
    _T_3177_im <= _T_3176_im;
    _T_3178_re <= _T_3177_re;
    _T_3178_im <= _T_3177_im;
    _T_3179_re <= _T_3178_re;
    _T_3179_im <= _T_3178_im;
    _T_3180_re <= _T_3179_re;
    _T_3180_im <= _T_3179_im;
    _T_3181_re <= _T_3180_re;
    _T_3181_im <= _T_3180_im;
    _T_3182_re <= _T_3181_re;
    _T_3182_im <= _T_3181_im;
    _T_3183_re <= _T_3182_re;
    _T_3183_im <= _T_3182_im;
    _T_3184_re <= _T_3183_re;
    _T_3184_im <= _T_3183_im;
    _T_3185_re <= _T_3184_re;
    _T_3185_im <= _T_3184_im;
    _T_3186_re <= _T_3185_re;
    _T_3186_im <= _T_3185_im;
    _T_3187_re <= _T_3186_re;
    _T_3187_im <= _T_3186_im;
    _T_3188_re <= _T_3187_re;
    _T_3188_im <= _T_3187_im;
    _T_3189_re <= _T_3188_re;
    _T_3189_im <= _T_3188_im;
    _T_3190_re <= _T_3189_re;
    _T_3190_im <= _T_3189_im;
    _T_3191_re <= _T_3190_re;
    _T_3191_im <= _T_3190_im;
    _T_3192_re <= _T_3191_re;
    _T_3192_im <= _T_3191_im;
    _T_3193_re <= _T_3192_re;
    _T_3193_im <= _T_3192_im;
    _T_3194_re <= _T_3193_re;
    _T_3194_im <= _T_3193_im;
    _T_3195_re <= _T_3194_re;
    _T_3195_im <= _T_3194_im;
    _T_3196_re <= _T_3195_re;
    _T_3196_im <= _T_3195_im;
    _T_3197_re <= _T_3196_re;
    _T_3197_im <= _T_3196_im;
    _T_3198_re <= _T_3197_re;
    _T_3198_im <= _T_3197_im;
    _T_3199_re <= _T_3198_re;
    _T_3199_im <= _T_3198_im;
    _T_3200_re <= _T_3199_re;
    _T_3200_im <= _T_3199_im;
    _T_3201_re <= _T_3200_re;
    _T_3201_im <= _T_3200_im;
    _T_3202_re <= _T_3201_re;
    _T_3202_im <= _T_3201_im;
    _T_3212_re <= Switch_4_io_out1_re;
    _T_3212_im <= Switch_4_io_out1_im;
    _T_3213_re <= _T_3212_re;
    _T_3213_im <= _T_3212_im;
    _T_3214_re <= _T_3213_re;
    _T_3214_im <= _T_3213_im;
    _T_3215_re <= _T_3214_re;
    _T_3215_im <= _T_3214_im;
    _T_3216_re <= _T_3215_re;
    _T_3216_im <= _T_3215_im;
    _T_3217_re <= _T_3216_re;
    _T_3217_im <= _T_3216_im;
    _T_3218_re <= _T_3217_re;
    _T_3218_im <= _T_3217_im;
    _T_3219_re <= _T_3218_re;
    _T_3219_im <= _T_3218_im;
    _T_3220_re <= _T_3219_re;
    _T_3220_im <= _T_3219_im;
    _T_3221_re <= _T_3220_re;
    _T_3221_im <= _T_3220_im;
    _T_3222_re <= _T_3221_re;
    _T_3222_im <= _T_3221_im;
    _T_3223_re <= _T_3222_re;
    _T_3223_im <= _T_3222_im;
    _T_3224_re <= _T_3223_re;
    _T_3224_im <= _T_3223_im;
    _T_3225_re <= _T_3224_re;
    _T_3225_im <= _T_3224_im;
    _T_3226_re <= _T_3225_re;
    _T_3226_im <= _T_3225_im;
    _T_3227_re <= _T_3226_re;
    _T_3227_im <= _T_3226_im;
    _T_3228_re <= _T_3227_re;
    _T_3228_im <= _T_3227_im;
    _T_3229_re <= _T_3228_re;
    _T_3229_im <= _T_3228_im;
    _T_3230_re <= _T_3229_re;
    _T_3230_im <= _T_3229_im;
    _T_3231_re <= _T_3230_re;
    _T_3231_im <= _T_3230_im;
    _T_3232_re <= _T_3231_re;
    _T_3232_im <= _T_3231_im;
    _T_3233_re <= _T_3232_re;
    _T_3233_im <= _T_3232_im;
    _T_3234_re <= _T_3233_re;
    _T_3234_im <= _T_3233_im;
    _T_3235_re <= _T_3234_re;
    _T_3235_im <= _T_3234_im;
    _T_3236_re <= _T_3235_re;
    _T_3236_im <= _T_3235_im;
    _T_3237_re <= _T_3236_re;
    _T_3237_im <= _T_3236_im;
    _T_3238_re <= _T_3237_re;
    _T_3238_im <= _T_3237_im;
    _T_3239_re <= _T_3238_re;
    _T_3239_im <= _T_3238_im;
    _T_3240_re <= _T_3239_re;
    _T_3240_im <= _T_3239_im;
    _T_3241_re <= _T_3240_re;
    _T_3241_im <= _T_3240_im;
    _T_3242_re <= _T_3241_re;
    _T_3242_im <= _T_3241_im;
    _T_3243_re <= _T_3242_re;
    _T_3243_im <= _T_3242_im;
    _T_3246_re <= Butterfly_5_io_out2_re;
    _T_3246_im <= Butterfly_5_io_out2_im;
    _T_3247_re <= _T_3246_re;
    _T_3247_im <= _T_3246_im;
    _T_3248_re <= _T_3247_re;
    _T_3248_im <= _T_3247_im;
    _T_3249_re <= _T_3248_re;
    _T_3249_im <= _T_3248_im;
    _T_3250_re <= _T_3249_re;
    _T_3250_im <= _T_3249_im;
    _T_3251_re <= _T_3250_re;
    _T_3251_im <= _T_3250_im;
    _T_3252_re <= _T_3251_re;
    _T_3252_im <= _T_3251_im;
    _T_3253_re <= _T_3252_re;
    _T_3253_im <= _T_3252_im;
    _T_3254_re <= _T_3253_re;
    _T_3254_im <= _T_3253_im;
    _T_3255_re <= _T_3254_re;
    _T_3255_im <= _T_3254_im;
    _T_3256_re <= _T_3255_re;
    _T_3256_im <= _T_3255_im;
    _T_3257_re <= _T_3256_re;
    _T_3257_im <= _T_3256_im;
    _T_3258_re <= _T_3257_re;
    _T_3258_im <= _T_3257_im;
    _T_3259_re <= _T_3258_re;
    _T_3259_im <= _T_3258_im;
    _T_3260_re <= _T_3259_re;
    _T_3260_im <= _T_3259_im;
    _T_3261_re <= _T_3260_re;
    _T_3261_im <= _T_3260_im;
    _T_3267_re <= Switch_5_io_out1_re;
    _T_3267_im <= Switch_5_io_out1_im;
    _T_3268_re <= _T_3267_re;
    _T_3268_im <= _T_3267_im;
    _T_3269_re <= _T_3268_re;
    _T_3269_im <= _T_3268_im;
    _T_3270_re <= _T_3269_re;
    _T_3270_im <= _T_3269_im;
    _T_3271_re <= _T_3270_re;
    _T_3271_im <= _T_3270_im;
    _T_3272_re <= _T_3271_re;
    _T_3272_im <= _T_3271_im;
    _T_3273_re <= _T_3272_re;
    _T_3273_im <= _T_3272_im;
    _T_3274_re <= _T_3273_re;
    _T_3274_im <= _T_3273_im;
    _T_3275_re <= _T_3274_re;
    _T_3275_im <= _T_3274_im;
    _T_3276_re <= _T_3275_re;
    _T_3276_im <= _T_3275_im;
    _T_3277_re <= _T_3276_re;
    _T_3277_im <= _T_3276_im;
    _T_3278_re <= _T_3277_re;
    _T_3278_im <= _T_3277_im;
    _T_3279_re <= _T_3278_re;
    _T_3279_im <= _T_3278_im;
    _T_3280_re <= _T_3279_re;
    _T_3280_im <= _T_3279_im;
    _T_3281_re <= _T_3280_re;
    _T_3281_im <= _T_3280_im;
    _T_3282_re <= _T_3281_re;
    _T_3282_im <= _T_3281_im;
    _T_3285_re <= Butterfly_6_io_out2_re;
    _T_3285_im <= Butterfly_6_io_out2_im;
    _T_3286_re <= _T_3285_re;
    _T_3286_im <= _T_3285_im;
    _T_3287_re <= _T_3286_re;
    _T_3287_im <= _T_3286_im;
    _T_3288_re <= _T_3287_re;
    _T_3288_im <= _T_3287_im;
    _T_3289_re <= _T_3288_re;
    _T_3289_im <= _T_3288_im;
    _T_3290_re <= _T_3289_re;
    _T_3290_im <= _T_3289_im;
    _T_3291_re <= _T_3290_re;
    _T_3291_im <= _T_3290_im;
    _T_3292_re <= _T_3291_re;
    _T_3292_im <= _T_3291_im;
    _T_3298_re <= Switch_6_io_out1_re;
    _T_3298_im <= Switch_6_io_out1_im;
    _T_3299_re <= _T_3298_re;
    _T_3299_im <= _T_3298_im;
    _T_3300_re <= _T_3299_re;
    _T_3300_im <= _T_3299_im;
    _T_3301_re <= _T_3300_re;
    _T_3301_im <= _T_3300_im;
    _T_3302_re <= _T_3301_re;
    _T_3302_im <= _T_3301_im;
    _T_3303_re <= _T_3302_re;
    _T_3303_im <= _T_3302_im;
    _T_3304_re <= _T_3303_re;
    _T_3304_im <= _T_3303_im;
    _T_3305_re <= _T_3304_re;
    _T_3305_im <= _T_3304_im;
    _T_3308_re <= Butterfly_7_io_out2_re;
    _T_3308_im <= Butterfly_7_io_out2_im;
    _T_3309_re <= _T_3308_re;
    _T_3309_im <= _T_3308_im;
    _T_3310_re <= _T_3309_re;
    _T_3310_im <= _T_3309_im;
    _T_3311_re <= _T_3310_re;
    _T_3311_im <= _T_3310_im;
    _T_3317_re <= Switch_7_io_out1_re;
    _T_3317_im <= Switch_7_io_out1_im;
    _T_3318_re <= _T_3317_re;
    _T_3318_im <= _T_3317_im;
    _T_3319_re <= _T_3318_re;
    _T_3319_im <= _T_3318_im;
    _T_3320_re <= _T_3319_re;
    _T_3320_im <= _T_3319_im;
    _T_3323_re <= Butterfly_8_io_out2_re;
    _T_3323_im <= Butterfly_8_io_out2_im;
    _T_3324_re <= _T_3323_re;
    _T_3324_im <= _T_3323_im;
    _T_3330_re <= Switch_8_io_out1_re;
    _T_3330_im <= Switch_8_io_out1_im;
    _T_3331_re <= _T_3330_re;
    _T_3331_im <= _T_3330_im;
    _T_3334_re <= Butterfly_9_io_out2_re;
    _T_3334_im <= Butterfly_9_io_out2_im;
    out1D1_re <= Switch_9_io_out1_re;
    out1D1_im <= Switch_9_io_out1_im;
    _T_3335_re <= ComplexAdd_io_res_re;
    _T_3335_im <= ComplexAdd_io_res_im;
    _T_3336_re <= ComplexSub_io_res_re;
    _T_3336_im <= ComplexSub_io_res_im;
  end
endmodule
