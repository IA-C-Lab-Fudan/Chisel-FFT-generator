module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T; // @[Butterfly.scala 57:28]
  wire [63:0] _T_1; // @[Butterfly.scala 57:52]
  wire [63:0] _T_4; // @[Butterfly.scala 57:40]
  wire [63:0] _T_5; // @[Butterfly.scala 58:28]
  wire [63:0] _T_6; // @[Butterfly.scala 58:52]
  wire [63:0] _T_9; // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2; // @[Butterfly.scala 58:15]
  assign _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  assign _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  assign _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  assign _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  assign _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  assign _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  assign _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT512RAM(
      input clk_in1_p,
    input clk_in1_n,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
    wire clock;
    clk_wiz_0 clk_wiz_0_inst0
       (
        // Clock out ports
        .clk_out1(clock),     // output clk_out1
       // Clock in ports
        .clk_in1_p(clk_in1_p),    // input clk_in1_p
        .clk_in1_n(clk_in1_n));    // input clk_in1_n
  wire  BRAM_clock; // @[FFT.scala 62:23]
  wire  BRAM_en; // @[FFT.scala 62:23]
  wire [7:0] BRAM_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_1_clock; // @[FFT.scala 62:23]
  wire  BRAM_1_en; // @[FFT.scala 62:23]
  wire [6:0] BRAM_1_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_1_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_2_clock; // @[FFT.scala 62:23]
  wire  BRAM_2_en; // @[FFT.scala 62:23]
  wire [5:0] BRAM_2_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_2_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire  BRAM_3_clock; // @[FFT.scala 62:23]
  wire  BRAM_3_en; // @[FFT.scala 62:23]
  wire [4:0] BRAM_3_addr; // @[FFT.scala 62:23]
  wire [63:0] BRAM_3_dout; // @[FFT.scala 62:23]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [8:0] cnt; // @[FFT.scala 40:20]
  reg [31:0] _RAND_0;
  wire [8:0] _T_1; // @[FFT.scala 42:16]
  reg [8:0] cntD1; // @[FFT.scala 44:22]
  reg [31:0] _RAND_1;
  reg [8:0] cntD2; // @[FFT.scala 45:22]
  reg [31:0] _RAND_2;
  reg [31:0] out1_0_re; // @[FFT.scala 50:23]
  reg [31:0] _RAND_3;
  reg [31:0] out1_0_im; // @[FFT.scala 50:23]
  reg [31:0] _RAND_4;
  reg [31:0] out2_0_re; // @[FFT.scala 51:23]
  reg [31:0] _RAND_5;
  reg [31:0] out2_0_im; // @[FFT.scala 51:23]
  reg [31:0] _RAND_6;
  wire [63:0] _T_148;
  reg [31:0] _T_153_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [31:0] _T_153_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [31:0] _T_154_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [31:0] _T_154_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [31:0] _T_155_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [31:0] _T_155_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg [31:0] _T_156_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg [31:0] _T_156_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg [31:0] _T_157_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] _T_157_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg [31:0] _T_158_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg [31:0] _T_158_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [31:0] _T_159_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] _T_159_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [31:0] _T_160_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] _T_160_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [31:0] _T_161_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [31:0] _T_162_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [31:0] _T_163_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg [31:0] _T_164_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg [31:0] _T_165_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg [31:0] _T_166_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [31:0] _T_167_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [31:0] _T_168_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [31:0] _T_169_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [31:0] _T_170_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [31:0] _T_171_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [31:0] _T_172_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg [31:0] _T_173_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] _T_174_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg [31:0] _T_175_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] _T_176_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] _T_177_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [31:0] _T_178_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [31:0] _T_179_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [31:0] _T_180_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg [31:0] _T_182_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg [31:0] _T_325_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg [31:0] _T_326_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg [31:0] _T_327_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg [31:0] _T_328_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_443;
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_444;
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_445;
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_446;
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_447;
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_448;
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_449;
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_450;
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_451;
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_452;
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_453;
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_454;
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_455;
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_456;
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_457;
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_458;
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_459;
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_460;
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_461;
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_462;
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_463;
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_464;
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_465;
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_466;
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_467;
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_468;
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_469;
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_470;
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_471;
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_472;
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_473;
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_474;
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_475;
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_476;
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_477;
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_478;
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_479;
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_480;
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_481;
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_482;
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_483;
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_484;
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_485;
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_486;
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_487;
  reg [31:0] _T_393_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_488;
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_489;
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_490;
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_491;
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_492;
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_493;
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_494;
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_495;
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_496;
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_497;
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_498;
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_499;
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_500;
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_501;
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_502;
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_503;
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_504;
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_505;
  reg [31:0] _T_402_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_506;
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_507;
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_508;
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_509;
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_510;
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_511;
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_512;
  reg [31:0] _T_406_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_513;
  reg [31:0] _T_406_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_514;
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_515;
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_516;
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_517;
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_518;
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_519;
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_520;
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_521;
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_522;
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_523;
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_524;
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_525;
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_526;
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_527;
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_528;
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_529;
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_530;
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_531;
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_532;
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_533;
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_534;
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_535;
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_536;
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_537;
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_538;
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_539;
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_540;
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_541;
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_542;
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_543;
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_544;
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_545;
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_546;
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_547;
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_548;
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_549;
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_550;
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_551;
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_552;
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_553;
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_554;
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_555;
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_556;
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_557;
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_558;
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_559;
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_560;
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_561;
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_562;
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_563;
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_564;
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_565;
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_566;
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_567;
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_568;
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_569;
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_570;
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_571;
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_572;
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_573;
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_574;
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_575;
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_576;
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_577;
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_578;
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_579;
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_580;
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_581;
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_582;
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_583;
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_584;
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_585;
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_586;
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_587;
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_588;
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_589;
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_590;
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_591;
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_592;
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_593;
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_594;
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_595;
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_596;
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_597;
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_598;
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_599;
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_600;
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_601;
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_602;
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_603;
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_604;
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_605;
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_606;
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_607;
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_608;
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_609;
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_610;
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_611;
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_612;
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_613;
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_614;
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_615;
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_616;
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_617;
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_618;
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_619;
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_620;
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_621;
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_622;
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_623;
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_624;
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_625;
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_626;
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_627;
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_628;
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_629;
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_630;
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_631;
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_632;
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_633;
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_634;
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_635;
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_636;
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_637;
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_638;
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_639;
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_640;
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_641;
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_642;
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_643;
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_644;
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_645;
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_646;
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_647;
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_648;
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_649;
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_650;
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_651;
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_652;
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_653;
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_654;
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_655;
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_656;
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_657;
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_658;
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_659;
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_660;
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_661;
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_662;
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_663;
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_664;
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_665;
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_666;
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_667;
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_668;
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_669;
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_670;
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_671;
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_672;
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_673;
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_674;
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_675;
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_676;
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_677;
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_678;
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_679;
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_680;
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_681;
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_682;
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_683;
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_684;
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_685;
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_686;
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_687;
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_688;
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_689;
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_690;
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_691;
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_692;
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_693;
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_694;
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_695;
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_696;
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_697;
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_698;
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_699;
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_700;
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_701;
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_702;
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_703;
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_704;
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_705;
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_706;
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_707;
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_708;
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_709;
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_710;
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_711;
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_712;
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_713;
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_714;
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_715;
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_716;
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_717;
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_718;
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_719;
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_720;
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_721;
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_722;
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_723;
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_724;
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_725;
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_726;
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_727;
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_728;
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_729;
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_730;
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_731;
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_732;
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_733;
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_734;
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_735;
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_736;
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_737;
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_738;
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_739;
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_740;
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_741;
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_742;
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_743;
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_744;
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_745;
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_746;
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_747;
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_748;
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_749;
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_750;
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_751;
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_752;
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_753;
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_754;
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_755;
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_756;
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_757;
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_758;
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_759;
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_760;
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_761;
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_762;
  reg [31:0] _T_533_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_763;
  reg [31:0] _T_533_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_764;
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_765;
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_766;
  reg [31:0] _T_535_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_767;
  reg [31:0] _T_535_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_768;
  reg [31:0] _T_536_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_769;
  reg [31:0] _T_536_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_770;
  reg [31:0] _T_537_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_771;
  reg [31:0] _T_537_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_772;
  reg [31:0] _T_538_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_773;
  reg [31:0] _T_538_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_774;
  wire [63:0] _T_543;
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_775;
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_776;
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_777;
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_778;
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_779;
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_780;
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_781;
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_782;
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_783;
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_784;
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_785;
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_786;
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_787;
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_788;
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_789;
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_790;
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_791;
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_792;
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_793;
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_794;
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_795;
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_796;
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_797;
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_798;
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_799;
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_800;
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_801;
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_802;
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_803;
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_804;
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_805;
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_806;
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_807;
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_808;
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_809;
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_810;
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_811;
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_812;
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_813;
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_814;
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_815;
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_816;
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_817;
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_818;
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_819;
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_820;
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_821;
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_822;
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_823;
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_824;
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_825;
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_826;
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_827;
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_828;
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_829;
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_830;
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_831;
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_832;
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_833;
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_834;
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_835;
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_836;
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_837;
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_838;
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_839;
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_840;
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_841;
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_842;
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_843;
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_844;
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_845;
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_846;
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_847;
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_848;
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_849;
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_850;
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_851;
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_852;
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_853;
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_854;
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_855;
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_856;
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_857;
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_858;
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_859;
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_860;
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_861;
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_862;
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_863;
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_864;
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_865;
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_866;
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_867;
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_868;
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_869;
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_870;
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_871;
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_872;
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_873;
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_874;
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_875;
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_876;
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_877;
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_878;
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_879;
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_880;
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_881;
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_882;
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_883;
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_884;
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_885;
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_886;
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_887;
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_888;
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_889;
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_890;
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_891;
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_892;
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_893;
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_894;
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_895;
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_896;
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_897;
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_898;
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_899;
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_900;
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_901;
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_902;
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_903;
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_904;
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_905;
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_906;
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_907;
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_908;
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_909;
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_910;
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_911;
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_912;
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_913;
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_914;
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_915;
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_916;
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_917;
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_918;
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_919;
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_920;
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_921;
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_922;
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_923;
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_924;
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_925;
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_926;
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_927;
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_928;
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_929;
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_930;
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_931;
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_932;
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_933;
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_934;
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_935;
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_936;
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_937;
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_938;
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_939;
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_940;
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_941;
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_942;
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_943;
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_944;
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_945;
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_946;
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_947;
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_948;
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_949;
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_950;
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_951;
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_952;
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_953;
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_954;
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_955;
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_956;
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_957;
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_958;
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_959;
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_960;
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_961;
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_962;
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_963;
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_964;
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_965;
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_966;
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_967;
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_968;
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_969;
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_970;
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_971;
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_972;
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_973;
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_974;
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_975;
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_976;
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_977;
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_978;
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_979;
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_980;
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_981;
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_982;
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_983;
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_984;
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_985;
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_986;
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_987;
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_988;
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_989;
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_990;
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_991;
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_992;
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_993;
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_994;
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_995;
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_996;
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_997;
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_998;
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_999;
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1000;
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1001;
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1002;
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1003;
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1004;
  reg [31:0] _T_663_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1005;
  reg [31:0] _T_663_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1006;
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1007;
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1008;
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1009;
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1010;
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1011;
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1012;
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1013;
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1014;
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1015;
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1016;
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1017;
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1018;
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1019;
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1020;
  reg [31:0] _T_671_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1021;
  reg [31:0] _T_671_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1022;
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1023;
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1024;
  reg [31:0] _T_673_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1025;
  reg [31:0] _T_673_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1026;
  reg [31:0] _T_674_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1027;
  reg [31:0] _T_674_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1028;
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1029;
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1030;
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1031;
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1032;
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1033;
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1034;
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1035;
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1036;
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1037;
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1038;
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1039;
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1040;
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1041;
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1042;
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1043;
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1044;
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1045;
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1046;
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1047;
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1048;
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1049;
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1050;
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1051;
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1052;
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1053;
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1054;
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1055;
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1056;
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1057;
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1058;
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1059;
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1060;
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1061;
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1062;
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1063;
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1064;
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1065;
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1066;
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1067;
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1068;
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1069;
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1070;
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1071;
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1072;
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1073;
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1074;
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1075;
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1076;
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1077;
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1078;
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1079;
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1080;
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1081;
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1082;
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1083;
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1084;
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1085;
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1086;
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1087;
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1088;
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1089;
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1090;
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1091;
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1092;
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1093;
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1094;
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1095;
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1096;
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1097;
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1098;
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1099;
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1100;
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1101;
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1102;
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1103;
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1104;
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1105;
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1106;
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1107;
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1108;
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1109;
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1110;
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1111;
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1112;
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1113;
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1114;
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1115;
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1116;
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1117;
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1118;
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1119;
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1120;
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1121;
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1122;
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1123;
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1124;
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1125;
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1126;
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1127;
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1128;
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1129;
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1130;
  reg [31:0] _T_728_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1131;
  reg [31:0] _T_728_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1132;
  reg [31:0] _T_729_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1133;
  reg [31:0] _T_729_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1134;
  reg [31:0] _T_730_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1135;
  reg [31:0] _T_730_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1136;
  reg [31:0] _T_731_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1137;
  reg [31:0] _T_731_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1138;
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1139;
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1140;
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1141;
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1142;
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1143;
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1144;
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1145;
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1146;
  reg [31:0] _T_736_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1147;
  reg [31:0] _T_736_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1148;
  reg [31:0] _T_737_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1149;
  reg [31:0] _T_737_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1150;
  reg [31:0] _T_738_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1151;
  reg [31:0] _T_738_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1152;
  reg [31:0] _T_739_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1153;
  reg [31:0] _T_739_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1154;
  reg [31:0] _T_740_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1155;
  reg [31:0] _T_740_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1156;
  reg [31:0] _T_741_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1157;
  reg [31:0] _T_741_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1158;
  wire [63:0] _T_746;
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1159;
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1160;
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1161;
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1162;
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1163;
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1164;
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1165;
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1166;
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1167;
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1168;
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1169;
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1170;
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1171;
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1172;
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1173;
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1174;
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1175;
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1176;
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1177;
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1178;
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1179;
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1180;
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1181;
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1182;
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1183;
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1184;
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1185;
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1186;
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1187;
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1188;
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1189;
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1190;
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1191;
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1192;
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1193;
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1194;
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1195;
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1196;
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1197;
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1198;
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1199;
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1200;
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1201;
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1202;
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1203;
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1204;
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1205;
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1206;
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1207;
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1208;
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1209;
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1210;
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1211;
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1212;
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1213;
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1214;
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1215;
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1216;
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1217;
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1218;
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1219;
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1220;
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1221;
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1222;
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1223;
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1224;
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1225;
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1226;
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1227;
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1228;
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1229;
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1230;
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1231;
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1232;
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1233;
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1234;
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1235;
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1236;
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1237;
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1238;
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1239;
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1240;
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1241;
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1242;
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1243;
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1244;
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1245;
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1246;
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1247;
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1248;
  reg [31:0] _T_796_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1249;
  reg [31:0] _T_796_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1250;
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1251;
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1252;
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1253;
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1254;
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1255;
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1256;
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1257;
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1258;
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1259;
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1260;
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1261;
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1262;
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1263;
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1264;
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1265;
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1266;
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1267;
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1268;
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1269;
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1270;
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1271;
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1272;
  reg [31:0] _T_808_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1273;
  reg [31:0] _T_808_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1274;
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1275;
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1276;
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1277;
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1278;
  reg [31:0] _T_811_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1279;
  reg [31:0] _T_811_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1280;
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1281;
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1282;
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1283;
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1284;
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1285;
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1286;
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1287;
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1288;
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1289;
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1290;
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1291;
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1292;
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1293;
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1294;
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1295;
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1296;
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1297;
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1298;
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1299;
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1300;
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1301;
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1302;
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1303;
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1304;
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1305;
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1306;
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1307;
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1308;
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1309;
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1310;
  reg [31:0] _T_829_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1311;
  reg [31:0] _T_829_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1312;
  reg [31:0] _T_830_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1313;
  reg [31:0] _T_830_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1314;
  reg [31:0] _T_831_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1315;
  reg [31:0] _T_831_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1316;
  reg [31:0] _T_832_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1317;
  reg [31:0] _T_832_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1318;
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1319;
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1320;
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1321;
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1322;
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1323;
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1324;
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1325;
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1326;
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1327;
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1328;
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1329;
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1330;
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1331;
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1332;
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1333;
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1334;
  reg [31:0] _T_841_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1335;
  reg [31:0] _T_841_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1336;
  reg [31:0] _T_842_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1337;
  reg [31:0] _T_842_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1338;
  reg [31:0] _T_843_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1339;
  reg [31:0] _T_843_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1340;
  reg [31:0] _T_844_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1341;
  reg [31:0] _T_844_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1342;
  reg [31:0] _T_845_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1343;
  reg [31:0] _T_845_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1344;
  reg [31:0] _T_846_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1345;
  reg [31:0] _T_846_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1346;
  reg [31:0] _T_847_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1347;
  reg [31:0] _T_847_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1348;
  reg [31:0] _T_848_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1349;
  reg [31:0] _T_848_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1350;
  wire [63:0] _T_853;
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1351;
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1352;
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1353;
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1354;
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1355;
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1356;
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1357;
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1358;
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1359;
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1360;
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1361;
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1362;
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1363;
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1364;
  reg [31:0] _T_865_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1365;
  reg [31:0] _T_865_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1366;
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1367;
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1368;
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1369;
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1370;
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1371;
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1372;
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1373;
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1374;
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1375;
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1376;
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1377;
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1378;
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1379;
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1380;
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1381;
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1382;
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1383;
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1384;
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1385;
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1386;
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1387;
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1388;
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1389;
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1390;
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1391;
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1392;
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1393;
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1394;
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1395;
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1396;
  reg [31:0] _T_881_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1397;
  reg [31:0] _T_881_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1398;
  reg [31:0] _T_882_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1399;
  reg [31:0] _T_882_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1400;
  reg [31:0] _T_883_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1401;
  reg [31:0] _T_883_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1402;
  reg [31:0] _T_884_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1403;
  reg [31:0] _T_884_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1404;
  reg [31:0] _T_885_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1405;
  reg [31:0] _T_885_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1406;
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1407;
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1408;
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1409;
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1410;
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1411;
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1412;
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1413;
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1414;
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1415;
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1416;
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1417;
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1418;
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1419;
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1420;
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1421;
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1422;
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1423;
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1424;
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1425;
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1426;
  reg [31:0] _T_898_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1427;
  reg [31:0] _T_898_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1428;
  reg [31:0] _T_899_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1429;
  reg [31:0] _T_899_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1430;
  reg [31:0] _T_900_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1431;
  reg [31:0] _T_900_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1432;
  reg [31:0] _T_901_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1433;
  reg [31:0] _T_901_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1434;
  reg [31:0] _T_902_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1435;
  reg [31:0] _T_902_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1436;
  reg [31:0] _T_903_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1437;
  reg [31:0] _T_903_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1438;
  reg [31:0] _T_904_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1439;
  reg [31:0] _T_904_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1440;
  reg [31:0] _T_905_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1441;
  reg [31:0] _T_905_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1442;
  reg [31:0] _T_906_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1443;
  reg [31:0] _T_906_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1444;
  reg [31:0] _T_907_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1445;
  reg [31:0] _T_907_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1446;
  wire [31:0] _GEN_1442; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1443; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1444; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1445; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1446; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1447; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1448; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1449; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1450; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1451; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1452; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1453; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1454; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1455; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1458; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1459; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1460; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1461; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1462; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1463; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1464; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1465; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1466; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1467; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1468; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1469; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1470; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1471; // @[FFT.scala 35:12]
  reg [31:0] _T_913_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1447;
  reg [31:0] _T_913_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1448;
  reg [31:0] _T_914_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1449;
  reg [31:0] _T_914_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1450;
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1451;
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1452;
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1453;
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1454;
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1455;
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1456;
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1457;
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1458;
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1459;
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1460;
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1461;
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1462;
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1463;
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1464;
  reg [31:0] _T_922_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1465;
  reg [31:0] _T_922_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1466;
  reg [31:0] _T_923_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1467;
  reg [31:0] _T_923_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1468;
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1469;
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1470;
  reg [31:0] _T_925_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1471;
  reg [31:0] _T_925_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1472;
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1473;
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1474;
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1475;
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1476;
  reg [31:0] _T_928_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1477;
  reg [31:0] _T_928_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1478;
  reg [31:0] _T_931_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1479;
  reg [31:0] _T_931_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1480;
  reg [31:0] _T_932_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1481;
  reg [31:0] _T_932_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1482;
  reg [31:0] _T_933_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1483;
  reg [31:0] _T_933_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1484;
  reg [31:0] _T_934_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1485;
  reg [31:0] _T_934_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1486;
  reg [31:0] _T_935_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1487;
  reg [31:0] _T_935_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1488;
  reg [31:0] _T_936_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1489;
  reg [31:0] _T_936_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1490;
  reg [31:0] _T_937_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1491;
  reg [31:0] _T_937_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1492;
  reg [31:0] _T_938_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1493;
  reg [31:0] _T_938_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1494;
  wire [31:0] _GEN_1522; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1523; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1524; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1525; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1526; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1527; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1530; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1531; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1532; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1533; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1534; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1535; // @[FFT.scala 35:12]
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1495;
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1496;
  reg [31:0] _T_945_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1497;
  reg [31:0] _T_945_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1498;
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1499;
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1500;
  reg [31:0] _T_947_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1501;
  reg [31:0] _T_947_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1502;
  reg [31:0] _T_948_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1503;
  reg [31:0] _T_948_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1504;
  reg [31:0] _T_949_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1505;
  reg [31:0] _T_949_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1506;
  reg [31:0] _T_950_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1507;
  reg [31:0] _T_950_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1508;
  reg [31:0] _T_951_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1509;
  reg [31:0] _T_951_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1510;
  reg [31:0] _T_954_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1511;
  reg [31:0] _T_954_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1512;
  reg [31:0] _T_955_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1513;
  reg [31:0] _T_955_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1514;
  reg [31:0] _T_956_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1515;
  reg [31:0] _T_956_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1516;
  reg [31:0] _T_957_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1517;
  reg [31:0] _T_957_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1518;
  wire [31:0] _GEN_1562; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1563; // @[FFT.scala 34:12]
  wire [31:0] _GEN_1566; // @[FFT.scala 35:12]
  wire [31:0] _GEN_1567; // @[FFT.scala 35:12]
  reg [31:0] _T_963_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1519;
  reg [31:0] _T_963_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1520;
  reg [31:0] _T_964_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1521;
  reg [31:0] _T_964_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1522;
  reg [31:0] _T_965_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1523;
  reg [31:0] _T_965_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1524;
  reg [31:0] _T_966_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1525;
  reg [31:0] _T_966_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1526;
  reg [31:0] _T_969_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1527;
  reg [31:0] _T_969_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1528;
  reg [31:0] _T_970_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1529;
  reg [31:0] _T_970_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1530;
  reg [31:0] _T_976_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1531;
  reg [31:0] _T_976_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1532;
  reg [31:0] _T_977_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1533;
  reg [31:0] _T_977_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1534;
  reg [31:0] _T_980_re; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1535;
  reg [31:0] _T_980_im; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1536;
  reg [31:0] out1D1_re; // @[FFT.scala 81:23]
  reg [31:0] _RAND_1537;
  reg [31:0] out1D1_im; // @[FFT.scala 81:23]
  reg [31:0] _RAND_1538;
  reg [31:0] _T_981_re; // @[FFT.scala 85:22]
  reg [31:0] _RAND_1539;
  reg [31:0] _T_981_im; // @[FFT.scala 85:22]
  reg [31:0] _RAND_1540;
  reg [31:0] _T_982_re; // @[FFT.scala 86:22]
  reg [31:0] _RAND_1541;
  reg [31:0] _T_982_im; // @[FFT.scala 86:22]
  reg [31:0] _RAND_1542;
  BRAM #(.ADDR_WIDTH(8), .DATA_WIDTH(64)) BRAM ( // @[FFT.scala 62:23]
    .clock(BRAM_clock),
    .en(BRAM_en),
    .addr(BRAM_addr),
    .dout(BRAM_dout)
  );
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(7), .DATA_WIDTH(64)) BRAM_1 ( // @[FFT.scala 62:23]
    .clock(BRAM_1_clock),
    .en(BRAM_1_en),
    .addr(BRAM_1_addr),
    .dout(BRAM_1_dout)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(6), .DATA_WIDTH(64)) BRAM_2 ( // @[FFT.scala 62:23]
    .clock(BRAM_2_clock),
    .en(BRAM_2_en),
    .addr(BRAM_2_addr),
    .dout(BRAM_2_dout)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  BRAM #(.ADDR_WIDTH(5), .DATA_WIDTH(64)) BRAM_3 ( // @[FFT.scala 62:23]
    .clock(BRAM_3_clock),
    .en(BRAM_3_en),
    .addr(BRAM_3_addr),
    .dout(BRAM_3_dout)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign _T_1 = cnt + 9'h1; // @[FFT.scala 42:16]
  assign _T_148 = BRAM_dout;
  assign _T_543 = BRAM_1_dout;
  assign _T_746 = BRAM_2_dout;
  assign _T_853 = BRAM_3_dout;
  assign _GEN_1442 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1443 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_1442); // @[FFT.scala 34:12]
  assign _GEN_1444 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_1443); // @[FFT.scala 34:12]
  assign _GEN_1445 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_1444); // @[FFT.scala 34:12]
  assign _GEN_1446 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_1445); // @[FFT.scala 34:12]
  assign _GEN_1447 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_1446); // @[FFT.scala 34:12]
  assign _GEN_1448 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_1447); // @[FFT.scala 34:12]
  assign _GEN_1449 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_1448); // @[FFT.scala 34:12]
  assign _GEN_1450 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_1449); // @[FFT.scala 34:12]
  assign _GEN_1451 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_1450); // @[FFT.scala 34:12]
  assign _GEN_1452 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1451); // @[FFT.scala 34:12]
  assign _GEN_1453 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_1452); // @[FFT.scala 34:12]
  assign _GEN_1454 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_1453); // @[FFT.scala 34:12]
  assign _GEN_1455 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_1454); // @[FFT.scala 34:12]
  assign _GEN_1458 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1459 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_1458); // @[FFT.scala 35:12]
  assign _GEN_1460 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1459); // @[FFT.scala 35:12]
  assign _GEN_1461 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_1460); // @[FFT.scala 35:12]
  assign _GEN_1462 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_1461); // @[FFT.scala 35:12]
  assign _GEN_1463 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_1462); // @[FFT.scala 35:12]
  assign _GEN_1464 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_1463); // @[FFT.scala 35:12]
  assign _GEN_1465 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_1464); // @[FFT.scala 35:12]
  assign _GEN_1466 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_1465); // @[FFT.scala 35:12]
  assign _GEN_1467 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_1466); // @[FFT.scala 35:12]
  assign _GEN_1468 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_1467); // @[FFT.scala 35:12]
  assign _GEN_1469 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_1468); // @[FFT.scala 35:12]
  assign _GEN_1470 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1469); // @[FFT.scala 35:12]
  assign _GEN_1471 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_1470); // @[FFT.scala 35:12]
  assign _GEN_1522 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1523 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_1522); // @[FFT.scala 34:12]
  assign _GEN_1524 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_1523); // @[FFT.scala 34:12]
  assign _GEN_1525 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_1524); // @[FFT.scala 34:12]
  assign _GEN_1526 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_1525); // @[FFT.scala 34:12]
  assign _GEN_1527 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_1526); // @[FFT.scala 34:12]
  assign _GEN_1530 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1531 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_1530); // @[FFT.scala 35:12]
  assign _GEN_1532 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_1531); // @[FFT.scala 35:12]
  assign _GEN_1533 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_1532); // @[FFT.scala 35:12]
  assign _GEN_1534 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_1533); // @[FFT.scala 35:12]
  assign _GEN_1535 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_1534); // @[FFT.scala 35:12]
  assign _GEN_1562 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 34:12]
  assign _GEN_1563 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_1562); // @[FFT.scala 34:12]
  assign _GEN_1566 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 35:12]
  assign _GEN_1567 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_1566); // @[FFT.scala 35:12]
  assign io_dOut1_re = _T_981_re; // @[FFT.scala 85:12]
  assign io_dOut1_im = _T_981_im; // @[FFT.scala 85:12]
  assign io_dOut2_re = _T_982_re; // @[FFT.scala 86:12]
  assign io_dOut2_im = _T_982_im; // @[FFT.scala 86:12]
  assign io_dout_valid = cntD2 == 9'h1ff; // @[FFT.scala 88:19]
  assign BRAM_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_addr = cnt[7:0]; // @[FFT.scala 64:19]
  assign Butterfly_io_in1_re = _T_408_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_408_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = out2_0_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = out2_0_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = _T_148[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = _T_148[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_538_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_538_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cntD1[7]; // @[Butterfly.scala 113:17]
  assign BRAM_1_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_1_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_1_addr = cnt[6:0]; // @[FFT.scala 64:19]
  assign Butterfly_1_io_in1_re = _T_675_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_675_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = _T_543[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = _T_543[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_741_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_741_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cntD1[6]; // @[Butterfly.scala 113:17]
  assign BRAM_2_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_2_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_2_addr = cnt[5:0]; // @[FFT.scala 64:19]
  assign Butterfly_2_io_in1_re = _T_814_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_814_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = _T_746[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = _T_746[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_848_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_848_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cntD1[5]; // @[Butterfly.scala 113:17]
  assign BRAM_3_clock = clock; // @[FFT.scala 65:20]
  assign BRAM_3_en = 1'h1; // @[FFT.scala 63:17]
  assign BRAM_3_addr = cnt[4:0]; // @[FFT.scala 64:19]
  assign Butterfly_3_io_in1_re = _T_889_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_889_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = _T_853[63:32]; // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = _T_853[31:0]; // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_907_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_907_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cntD1[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_928_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_928_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_1455); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_1471); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_938_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_938_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cntD1[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_951_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_951_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_1527); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_1535); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_957_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_957_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cntD1[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_966_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_966_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_1563); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_1567); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_970_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_970_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cntD1[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_7_io_in1_re = _T_977_re; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in1_im = _T_977_im; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_7_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in2_re = _T_980_re; // @[Butterfly.scala 112:17]
  assign Switch_7_io_in2_im = _T_980_im; // @[Butterfly.scala 112:17]
  assign Switch_7_io_sel = cntD1[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntD1 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cntD2 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out1_0_re = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out1_0_im = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out2_0_re = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out2_0_im = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_153_re = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_153_im = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_154_re = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_154_im = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_155_re = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_155_im = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_156_re = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_156_im = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_157_re = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_157_im = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_158_re = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_158_im = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_159_re = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_159_im = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_160_re = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_160_im = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_161_re = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_161_im = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_162_re = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_162_im = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_163_re = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_163_im = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_164_re = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_164_im = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_165_re = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_165_im = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_166_re = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_166_im = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_167_re = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_167_im = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_168_re = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_168_im = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_169_re = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_169_im = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_170_re = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_170_im = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_171_re = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_171_im = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_172_re = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_172_im = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_173_re = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_173_im = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_174_re = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_174_im = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_175_re = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_175_im = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_176_re = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_176_im = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_177_re = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_177_im = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_178_re = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_178_im = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_179_re = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_179_im = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_180_re = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_180_im = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_181_re = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_181_im = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_182_re = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_182_im = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_183_re = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_183_im = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_184_re = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_184_im = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_185_re = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_185_im = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_186_re = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_186_im = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_187_re = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_187_im = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_188_re = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_188_im = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_189_re = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_189_im = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_190_re = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_190_im = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_191_re = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_191_im = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_192_re = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_192_im = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_193_re = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_193_im = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_194_re = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_194_im = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_195_re = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_195_im = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_196_re = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_196_im = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_197_re = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_197_im = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_198_re = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_198_im = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_199_re = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_199_im = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_200_re = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_200_im = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_201_re = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_201_im = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_202_re = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_202_im = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_203_re = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_203_im = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_204_re = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_204_im = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_205_re = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_205_im = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_206_re = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_206_im = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_207_re = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_207_im = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_208_re = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_208_im = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_209_re = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_209_im = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_210_re = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_210_im = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_211_re = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_211_im = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_212_re = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_212_im = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_213_re = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_213_im = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_214_re = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_214_im = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_215_re = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_215_im = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_216_re = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_216_im = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_217_re = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_217_im = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_218_re = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_218_im = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_219_re = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_219_im = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_220_re = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_220_im = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_221_re = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_221_im = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_222_re = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_222_im = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_223_re = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_223_im = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_224_re = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_224_im = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_225_re = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_225_im = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_226_re = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_226_im = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_227_re = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_227_im = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_228_re = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_228_im = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_229_re = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_229_im = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_230_re = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_230_im = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_231_re = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_231_im = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_232_re = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_232_im = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_233_re = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_233_im = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_234_re = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_234_im = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_235_re = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_235_im = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_236_re = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_236_im = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_237_re = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_237_im = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_238_re = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_238_im = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_239_re = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_239_im = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_240_re = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_240_im = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_241_re = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_241_im = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_242_re = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_242_im = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_243_re = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_243_im = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_244_re = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_244_im = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_245_re = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_245_im = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_246_re = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_246_im = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_247_re = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_247_im = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_248_re = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_248_im = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_249_re = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_249_im = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_250_re = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_250_im = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_251_re = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_251_im = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_252_re = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_252_im = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_253_re = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_253_im = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_254_re = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_254_im = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_255_re = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_255_im = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_256_re = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_256_im = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_257_re = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_257_im = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_258_re = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_258_im = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_259_re = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_259_im = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_260_re = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_260_im = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_261_re = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_261_im = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_262_re = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_262_im = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_263_re = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_263_im = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_264_re = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_264_im = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_265_re = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_265_im = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_266_re = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_266_im = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_267_re = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_267_im = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_268_re = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_268_im = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_269_re = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_269_im = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_270_re = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_270_im = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_271_re = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_271_im = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_272_re = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_272_im = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_273_re = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_273_im = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_274_re = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_274_im = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_275_re = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_275_im = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_276_re = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_276_im = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_277_re = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_277_im = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_278_re = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_278_im = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_279_re = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_279_im = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_280_re = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_280_im = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_281_re = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_281_im = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_282_re = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_282_im = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_283_re = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_283_im = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_284_re = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_284_im = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_285_re = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_285_im = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_286_re = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_286_im = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_287_re = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_287_im = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_288_re = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_288_im = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_289_re = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_289_im = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_290_re = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_290_im = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_291_re = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_291_im = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_292_re = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_292_im = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_293_re = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_293_im = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_294_re = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_294_im = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_295_re = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_295_im = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_296_re = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_296_im = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_297_re = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_297_im = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_298_re = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_298_im = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_299_re = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_299_im = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_300_re = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_300_im = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_301_re = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_301_im = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_302_re = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_302_im = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_303_re = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_303_im = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_304_re = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_304_im = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_305_re = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_305_im = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_306_re = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_306_im = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_307_re = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_307_im = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_308_re = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_308_im = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_309_re = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_309_im = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_310_re = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_310_im = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_311_re = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_311_im = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_312_re = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_312_im = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_313_re = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_313_im = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_314_re = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_314_im = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_315_re = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_315_im = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_316_re = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_316_im = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_317_re = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_317_im = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_318_re = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_318_im = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_319_re = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_319_im = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_320_re = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_320_im = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_321_re = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_321_im = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_322_re = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_322_im = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_323_re = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_323_im = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_324_re = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_324_im = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_325_re = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_325_im = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_326_re = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_326_im = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_327_re = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_327_im = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_328_re = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_328_im = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_329_re = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_329_im = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_330_re = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_330_im = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_331_re = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_331_im = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_332_re = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_332_im = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_333_re = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_333_im = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_334_re = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_334_im = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_335_re = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_335_im = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_336_re = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_336_im = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_337_re = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_337_im = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_338_re = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_338_im = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_339_re = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_339_im = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_340_re = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_340_im = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_341_re = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_341_im = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_342_re = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_342_im = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_343_re = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_343_im = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_344_re = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_344_im = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_345_re = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_345_im = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_346_re = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_346_im = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_347_re = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_347_im = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_348_re = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_348_im = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_349_re = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_349_im = _RAND_400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_350_re = _RAND_401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_350_im = _RAND_402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_351_re = _RAND_403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_351_im = _RAND_404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_352_re = _RAND_405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_352_im = _RAND_406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_353_re = _RAND_407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_353_im = _RAND_408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_354_re = _RAND_409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_354_im = _RAND_410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_355_re = _RAND_411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_355_im = _RAND_412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_356_re = _RAND_413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_356_im = _RAND_414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_357_re = _RAND_415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_357_im = _RAND_416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_358_re = _RAND_417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_358_im = _RAND_418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_359_re = _RAND_419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_359_im = _RAND_420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_360_re = _RAND_421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_360_im = _RAND_422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_361_re = _RAND_423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_361_im = _RAND_424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_362_re = _RAND_425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_362_im = _RAND_426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_363_re = _RAND_427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_363_im = _RAND_428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_364_re = _RAND_429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_364_im = _RAND_430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_365_re = _RAND_431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_365_im = _RAND_432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_366_re = _RAND_433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_366_im = _RAND_434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_367_re = _RAND_435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_367_im = _RAND_436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_368_re = _RAND_437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_368_im = _RAND_438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_369_re = _RAND_439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_369_im = _RAND_440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_370_re = _RAND_441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_370_im = _RAND_442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_371_re = _RAND_443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_371_im = _RAND_444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_372_re = _RAND_445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_372_im = _RAND_446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_373_re = _RAND_447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_373_im = _RAND_448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_374_re = _RAND_449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_374_im = _RAND_450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_375_re = _RAND_451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_375_im = _RAND_452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_376_re = _RAND_453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_376_im = _RAND_454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_377_re = _RAND_455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_377_im = _RAND_456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_378_re = _RAND_457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_378_im = _RAND_458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_379_re = _RAND_459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_379_im = _RAND_460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_380_re = _RAND_461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_380_im = _RAND_462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_381_re = _RAND_463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_381_im = _RAND_464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_382_re = _RAND_465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_382_im = _RAND_466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_383_re = _RAND_467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_383_im = _RAND_468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_384_re = _RAND_469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_384_im = _RAND_470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_385_re = _RAND_471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_385_im = _RAND_472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_386_re = _RAND_473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_386_im = _RAND_474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_387_re = _RAND_475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_387_im = _RAND_476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_388_re = _RAND_477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_388_im = _RAND_478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_389_re = _RAND_479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_389_im = _RAND_480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_390_re = _RAND_481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_390_im = _RAND_482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_391_re = _RAND_483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_391_im = _RAND_484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_392_re = _RAND_485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_392_im = _RAND_486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_393_re = _RAND_487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_393_im = _RAND_488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_394_re = _RAND_489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_394_im = _RAND_490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_395_re = _RAND_491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_395_im = _RAND_492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_396_re = _RAND_493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_396_im = _RAND_494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_397_re = _RAND_495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_397_im = _RAND_496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_398_re = _RAND_497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_398_im = _RAND_498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_399_re = _RAND_499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_399_im = _RAND_500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_400_re = _RAND_501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_400_im = _RAND_502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_401_re = _RAND_503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_401_im = _RAND_504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_402_re = _RAND_505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_402_im = _RAND_506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_403_re = _RAND_507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_403_im = _RAND_508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_404_re = _RAND_509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_404_im = _RAND_510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_405_re = _RAND_511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_405_im = _RAND_512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_406_re = _RAND_513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_406_im = _RAND_514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_407_re = _RAND_515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_407_im = _RAND_516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_408_re = _RAND_517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_408_im = _RAND_518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_411_re = _RAND_519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_411_im = _RAND_520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_412_re = _RAND_521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_412_im = _RAND_522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_413_re = _RAND_523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_413_im = _RAND_524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_414_re = _RAND_525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_414_im = _RAND_526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_415_re = _RAND_527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_415_im = _RAND_528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_416_re = _RAND_529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_416_im = _RAND_530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_417_re = _RAND_531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_417_im = _RAND_532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_418_re = _RAND_533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_418_im = _RAND_534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_419_re = _RAND_535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_419_im = _RAND_536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_420_re = _RAND_537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_420_im = _RAND_538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_421_re = _RAND_539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_421_im = _RAND_540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_422_re = _RAND_541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_422_im = _RAND_542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_423_re = _RAND_543[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_423_im = _RAND_544[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_424_re = _RAND_545[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_424_im = _RAND_546[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_425_re = _RAND_547[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_425_im = _RAND_548[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_426_re = _RAND_549[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_426_im = _RAND_550[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_427_re = _RAND_551[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_427_im = _RAND_552[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_428_re = _RAND_553[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_428_im = _RAND_554[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_429_re = _RAND_555[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_429_im = _RAND_556[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_430_re = _RAND_557[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_430_im = _RAND_558[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_431_re = _RAND_559[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_431_im = _RAND_560[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_432_re = _RAND_561[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_432_im = _RAND_562[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_433_re = _RAND_563[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_433_im = _RAND_564[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_434_re = _RAND_565[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_434_im = _RAND_566[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_435_re = _RAND_567[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_435_im = _RAND_568[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_436_re = _RAND_569[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_436_im = _RAND_570[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_437_re = _RAND_571[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_437_im = _RAND_572[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_438_re = _RAND_573[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_438_im = _RAND_574[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_439_re = _RAND_575[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_439_im = _RAND_576[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_440_re = _RAND_577[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_440_im = _RAND_578[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_441_re = _RAND_579[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_441_im = _RAND_580[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_442_re = _RAND_581[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_442_im = _RAND_582[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_443_re = _RAND_583[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_443_im = _RAND_584[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_444_re = _RAND_585[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_444_im = _RAND_586[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_445_re = _RAND_587[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_445_im = _RAND_588[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_446_re = _RAND_589[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_446_im = _RAND_590[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_447_re = _RAND_591[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_447_im = _RAND_592[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_448_re = _RAND_593[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_448_im = _RAND_594[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_449_re = _RAND_595[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_449_im = _RAND_596[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_450_re = _RAND_597[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_450_im = _RAND_598[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_451_re = _RAND_599[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_451_im = _RAND_600[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_452_re = _RAND_601[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_452_im = _RAND_602[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_453_re = _RAND_603[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_453_im = _RAND_604[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_454_re = _RAND_605[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_454_im = _RAND_606[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_455_re = _RAND_607[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_455_im = _RAND_608[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_456_re = _RAND_609[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_456_im = _RAND_610[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_457_re = _RAND_611[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_457_im = _RAND_612[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_458_re = _RAND_613[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_458_im = _RAND_614[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_459_re = _RAND_615[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_459_im = _RAND_616[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_460_re = _RAND_617[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_460_im = _RAND_618[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_461_re = _RAND_619[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_461_im = _RAND_620[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_462_re = _RAND_621[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_462_im = _RAND_622[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_463_re = _RAND_623[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_463_im = _RAND_624[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_464_re = _RAND_625[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_464_im = _RAND_626[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_465_re = _RAND_627[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_465_im = _RAND_628[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_466_re = _RAND_629[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_466_im = _RAND_630[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_467_re = _RAND_631[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_467_im = _RAND_632[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_468_re = _RAND_633[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_468_im = _RAND_634[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_469_re = _RAND_635[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_469_im = _RAND_636[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_470_re = _RAND_637[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_470_im = _RAND_638[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_471_re = _RAND_639[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_471_im = _RAND_640[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_472_re = _RAND_641[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_472_im = _RAND_642[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_473_re = _RAND_643[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_473_im = _RAND_644[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_474_re = _RAND_645[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_474_im = _RAND_646[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_475_re = _RAND_647[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_475_im = _RAND_648[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_476_re = _RAND_649[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_476_im = _RAND_650[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_477_re = _RAND_651[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_477_im = _RAND_652[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_478_re = _RAND_653[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_478_im = _RAND_654[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_479_re = _RAND_655[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_479_im = _RAND_656[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_480_re = _RAND_657[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_480_im = _RAND_658[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_481_re = _RAND_659[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_481_im = _RAND_660[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_482_re = _RAND_661[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_482_im = _RAND_662[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_483_re = _RAND_663[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_483_im = _RAND_664[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_484_re = _RAND_665[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_484_im = _RAND_666[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_485_re = _RAND_667[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_485_im = _RAND_668[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_486_re = _RAND_669[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_486_im = _RAND_670[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_487_re = _RAND_671[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_487_im = _RAND_672[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_488_re = _RAND_673[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_488_im = _RAND_674[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_489_re = _RAND_675[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_489_im = _RAND_676[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_490_re = _RAND_677[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_490_im = _RAND_678[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_491_re = _RAND_679[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_491_im = _RAND_680[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_492_re = _RAND_681[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_492_im = _RAND_682[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_493_re = _RAND_683[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_493_im = _RAND_684[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_494_re = _RAND_685[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_494_im = _RAND_686[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_495_re = _RAND_687[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_495_im = _RAND_688[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_496_re = _RAND_689[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_496_im = _RAND_690[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_497_re = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_497_im = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_498_re = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_498_im = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_499_re = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_499_im = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_500_re = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_500_im = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_501_re = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_501_im = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_502_re = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_502_im = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_503_re = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_503_im = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_504_re = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_504_im = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_505_re = _RAND_707[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_505_im = _RAND_708[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_506_re = _RAND_709[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_506_im = _RAND_710[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_507_re = _RAND_711[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_507_im = _RAND_712[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_508_re = _RAND_713[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_508_im = _RAND_714[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_509_re = _RAND_715[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_509_im = _RAND_716[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_510_re = _RAND_717[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_510_im = _RAND_718[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_511_re = _RAND_719[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_511_im = _RAND_720[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_512_re = _RAND_721[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_512_im = _RAND_722[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_513_re = _RAND_723[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_513_im = _RAND_724[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_514_re = _RAND_725[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_514_im = _RAND_726[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_515_re = _RAND_727[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_515_im = _RAND_728[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_516_re = _RAND_729[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_516_im = _RAND_730[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_517_re = _RAND_731[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_517_im = _RAND_732[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_518_re = _RAND_733[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_518_im = _RAND_734[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_519_re = _RAND_735[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_519_im = _RAND_736[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_520_re = _RAND_737[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_520_im = _RAND_738[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_521_re = _RAND_739[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_521_im = _RAND_740[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_522_re = _RAND_741[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_522_im = _RAND_742[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_523_re = _RAND_743[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_523_im = _RAND_744[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_524_re = _RAND_745[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_524_im = _RAND_746[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_525_re = _RAND_747[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_525_im = _RAND_748[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_526_re = _RAND_749[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_526_im = _RAND_750[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_527_re = _RAND_751[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_527_im = _RAND_752[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_528_re = _RAND_753[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_528_im = _RAND_754[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_529_re = _RAND_755[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_529_im = _RAND_756[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_530_re = _RAND_757[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_530_im = _RAND_758[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_531_re = _RAND_759[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_531_im = _RAND_760[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_532_re = _RAND_761[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_532_im = _RAND_762[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_533_re = _RAND_763[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_533_im = _RAND_764[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_534_re = _RAND_765[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_534_im = _RAND_766[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_535_re = _RAND_767[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_535_im = _RAND_768[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_536_re = _RAND_769[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_536_im = _RAND_770[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_537_re = _RAND_771[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_537_im = _RAND_772[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_538_re = _RAND_773[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_538_im = _RAND_774[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_548_re = _RAND_775[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_548_im = _RAND_776[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_549_re = _RAND_777[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_549_im = _RAND_778[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_550_re = _RAND_779[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_550_im = _RAND_780[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_551_re = _RAND_781[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_551_im = _RAND_782[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_552_re = _RAND_783[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_552_im = _RAND_784[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_553_re = _RAND_785[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_553_im = _RAND_786[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_554_re = _RAND_787[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_554_im = _RAND_788[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_555_re = _RAND_789[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_555_im = _RAND_790[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_556_re = _RAND_791[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_556_im = _RAND_792[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_557_re = _RAND_793[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_557_im = _RAND_794[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_558_re = _RAND_795[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_558_im = _RAND_796[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_559_re = _RAND_797[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_559_im = _RAND_798[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_560_re = _RAND_799[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_560_im = _RAND_800[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_561_re = _RAND_801[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_561_im = _RAND_802[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_562_re = _RAND_803[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_562_im = _RAND_804[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_563_re = _RAND_805[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_563_im = _RAND_806[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_564_re = _RAND_807[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_564_im = _RAND_808[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_565_re = _RAND_809[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_565_im = _RAND_810[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_566_re = _RAND_811[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_566_im = _RAND_812[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_567_re = _RAND_813[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_567_im = _RAND_814[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_568_re = _RAND_815[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_568_im = _RAND_816[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_569_re = _RAND_817[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_569_im = _RAND_818[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_570_re = _RAND_819[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_570_im = _RAND_820[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_571_re = _RAND_821[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_571_im = _RAND_822[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_572_re = _RAND_823[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_572_im = _RAND_824[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_573_re = _RAND_825[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_573_im = _RAND_826[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_574_re = _RAND_827[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_574_im = _RAND_828[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_575_re = _RAND_829[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_575_im = _RAND_830[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_576_re = _RAND_831[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_576_im = _RAND_832[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_577_re = _RAND_833[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_577_im = _RAND_834[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_578_re = _RAND_835[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_578_im = _RAND_836[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_579_re = _RAND_837[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_579_im = _RAND_838[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_580_re = _RAND_839[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_580_im = _RAND_840[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_581_re = _RAND_841[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_581_im = _RAND_842[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_582_re = _RAND_843[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_582_im = _RAND_844[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_583_re = _RAND_845[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_583_im = _RAND_846[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_584_re = _RAND_847[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_584_im = _RAND_848[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_585_re = _RAND_849[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_585_im = _RAND_850[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_586_re = _RAND_851[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_586_im = _RAND_852[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_587_re = _RAND_853[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_587_im = _RAND_854[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_588_re = _RAND_855[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_588_im = _RAND_856[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_589_re = _RAND_857[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_589_im = _RAND_858[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_590_re = _RAND_859[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_590_im = _RAND_860[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_591_re = _RAND_861[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_591_im = _RAND_862[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_592_re = _RAND_863[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_592_im = _RAND_864[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_593_re = _RAND_865[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_593_im = _RAND_866[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_594_re = _RAND_867[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_594_im = _RAND_868[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_595_re = _RAND_869[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_595_im = _RAND_870[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_596_re = _RAND_871[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_596_im = _RAND_872[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_597_re = _RAND_873[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_597_im = _RAND_874[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_598_re = _RAND_875[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_598_im = _RAND_876[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_599_re = _RAND_877[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_599_im = _RAND_878[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_600_re = _RAND_879[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_600_im = _RAND_880[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_601_re = _RAND_881[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_601_im = _RAND_882[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_602_re = _RAND_883[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_602_im = _RAND_884[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_603_re = _RAND_885[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_603_im = _RAND_886[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_604_re = _RAND_887[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_604_im = _RAND_888[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_605_re = _RAND_889[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_605_im = _RAND_890[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_606_re = _RAND_891[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_606_im = _RAND_892[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_607_re = _RAND_893[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_607_im = _RAND_894[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_608_re = _RAND_895[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_608_im = _RAND_896[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_609_re = _RAND_897[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_609_im = _RAND_898[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_610_re = _RAND_899[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_610_im = _RAND_900[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_611_re = _RAND_901[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_611_im = _RAND_902[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_612_re = _RAND_903[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_612_im = _RAND_904[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_613_re = _RAND_905[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_613_im = _RAND_906[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_614_re = _RAND_907[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_614_im = _RAND_908[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_615_re = _RAND_909[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_615_im = _RAND_910[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_616_re = _RAND_911[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_616_im = _RAND_912[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_617_re = _RAND_913[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_617_im = _RAND_914[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_618_re = _RAND_915[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_618_im = _RAND_916[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_619_re = _RAND_917[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_619_im = _RAND_918[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_620_re = _RAND_919[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_620_im = _RAND_920[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_621_re = _RAND_921[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_621_im = _RAND_922[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_622_re = _RAND_923[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_622_im = _RAND_924[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_623_re = _RAND_925[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_623_im = _RAND_926[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_624_re = _RAND_927[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_624_im = _RAND_928[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_625_re = _RAND_929[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_625_im = _RAND_930[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_626_re = _RAND_931[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_626_im = _RAND_932[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_627_re = _RAND_933[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_627_im = _RAND_934[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_628_re = _RAND_935[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_628_im = _RAND_936[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_629_re = _RAND_937[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_629_im = _RAND_938[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_630_re = _RAND_939[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_630_im = _RAND_940[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_631_re = _RAND_941[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_631_im = _RAND_942[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_632_re = _RAND_943[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_632_im = _RAND_944[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_633_re = _RAND_945[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_633_im = _RAND_946[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_634_re = _RAND_947[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_634_im = _RAND_948[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_635_re = _RAND_949[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_635_im = _RAND_950[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_636_re = _RAND_951[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_636_im = _RAND_952[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_637_re = _RAND_953[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_637_im = _RAND_954[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_638_re = _RAND_955[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_638_im = _RAND_956[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_639_re = _RAND_957[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_639_im = _RAND_958[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_640_re = _RAND_959[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_640_im = _RAND_960[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_641_re = _RAND_961[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_641_im = _RAND_962[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_642_re = _RAND_963[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_642_im = _RAND_964[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_643_re = _RAND_965[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_643_im = _RAND_966[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_644_re = _RAND_967[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_644_im = _RAND_968[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_645_re = _RAND_969[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_645_im = _RAND_970[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_646_re = _RAND_971[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_646_im = _RAND_972[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_647_re = _RAND_973[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_647_im = _RAND_974[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_648_re = _RAND_975[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_648_im = _RAND_976[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_649_re = _RAND_977[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_649_im = _RAND_978[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_650_re = _RAND_979[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_650_im = _RAND_980[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_651_re = _RAND_981[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_651_im = _RAND_982[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_652_re = _RAND_983[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_652_im = _RAND_984[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_653_re = _RAND_985[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_653_im = _RAND_986[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_654_re = _RAND_987[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_654_im = _RAND_988[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_655_re = _RAND_989[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_655_im = _RAND_990[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_656_re = _RAND_991[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_656_im = _RAND_992[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_657_re = _RAND_993[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_657_im = _RAND_994[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_658_re = _RAND_995[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_658_im = _RAND_996[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_659_re = _RAND_997[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_659_im = _RAND_998[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_660_re = _RAND_999[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_660_im = _RAND_1000[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_661_re = _RAND_1001[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_661_im = _RAND_1002[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_662_re = _RAND_1003[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_662_im = _RAND_1004[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_663_re = _RAND_1005[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_663_im = _RAND_1006[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_664_re = _RAND_1007[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_664_im = _RAND_1008[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_665_re = _RAND_1009[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_665_im = _RAND_1010[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_666_re = _RAND_1011[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_666_im = _RAND_1012[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_667_re = _RAND_1013[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_667_im = _RAND_1014[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_668_re = _RAND_1015[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_668_im = _RAND_1016[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_669_re = _RAND_1017[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_669_im = _RAND_1018[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_670_re = _RAND_1019[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_670_im = _RAND_1020[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_671_re = _RAND_1021[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_671_im = _RAND_1022[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_672_re = _RAND_1023[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_672_im = _RAND_1024[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_673_re = _RAND_1025[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_673_im = _RAND_1026[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_674_re = _RAND_1027[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_674_im = _RAND_1028[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_675_re = _RAND_1029[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_675_im = _RAND_1030[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_678_re = _RAND_1031[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_678_im = _RAND_1032[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_679_re = _RAND_1033[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_679_im = _RAND_1034[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_680_re = _RAND_1035[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_680_im = _RAND_1036[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_681_re = _RAND_1037[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_681_im = _RAND_1038[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_682_re = _RAND_1039[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_682_im = _RAND_1040[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_683_re = _RAND_1041[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_683_im = _RAND_1042[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_684_re = _RAND_1043[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_684_im = _RAND_1044[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_685_re = _RAND_1045[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_685_im = _RAND_1046[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_686_re = _RAND_1047[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_686_im = _RAND_1048[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_687_re = _RAND_1049[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_687_im = _RAND_1050[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_688_re = _RAND_1051[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_688_im = _RAND_1052[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_689_re = _RAND_1053[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_689_im = _RAND_1054[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_690_re = _RAND_1055[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_690_im = _RAND_1056[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_691_re = _RAND_1057[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_691_im = _RAND_1058[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_692_re = _RAND_1059[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_692_im = _RAND_1060[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_693_re = _RAND_1061[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_693_im = _RAND_1062[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_694_re = _RAND_1063[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_694_im = _RAND_1064[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_695_re = _RAND_1065[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_695_im = _RAND_1066[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_696_re = _RAND_1067[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_696_im = _RAND_1068[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_697_re = _RAND_1069[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_697_im = _RAND_1070[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_698_re = _RAND_1071[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_698_im = _RAND_1072[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_699_re = _RAND_1073[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_699_im = _RAND_1074[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_700_re = _RAND_1075[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_700_im = _RAND_1076[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_701_re = _RAND_1077[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_701_im = _RAND_1078[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_702_re = _RAND_1079[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_702_im = _RAND_1080[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_703_re = _RAND_1081[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_703_im = _RAND_1082[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_704_re = _RAND_1083[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_704_im = _RAND_1084[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_705_re = _RAND_1085[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_705_im = _RAND_1086[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_706_re = _RAND_1087[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_706_im = _RAND_1088[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_707_re = _RAND_1089[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_707_im = _RAND_1090[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_708_re = _RAND_1091[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_708_im = _RAND_1092[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_709_re = _RAND_1093[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_709_im = _RAND_1094[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_710_re = _RAND_1095[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_710_im = _RAND_1096[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_711_re = _RAND_1097[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_711_im = _RAND_1098[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_712_re = _RAND_1099[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_712_im = _RAND_1100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_713_re = _RAND_1101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_713_im = _RAND_1102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_714_re = _RAND_1103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_714_im = _RAND_1104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_715_re = _RAND_1105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_715_im = _RAND_1106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_716_re = _RAND_1107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_716_im = _RAND_1108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_717_re = _RAND_1109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_717_im = _RAND_1110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_718_re = _RAND_1111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_718_im = _RAND_1112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_719_re = _RAND_1113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_719_im = _RAND_1114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_720_re = _RAND_1115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_720_im = _RAND_1116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_721_re = _RAND_1117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_721_im = _RAND_1118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_722_re = _RAND_1119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_722_im = _RAND_1120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_723_re = _RAND_1121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_723_im = _RAND_1122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_724_re = _RAND_1123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_724_im = _RAND_1124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_725_re = _RAND_1125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_725_im = _RAND_1126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_726_re = _RAND_1127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_726_im = _RAND_1128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_727_re = _RAND_1129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_727_im = _RAND_1130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_728_re = _RAND_1131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_728_im = _RAND_1132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_729_re = _RAND_1133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_729_im = _RAND_1134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_730_re = _RAND_1135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_730_im = _RAND_1136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_731_re = _RAND_1137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_731_im = _RAND_1138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_732_re = _RAND_1139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_732_im = _RAND_1140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_733_re = _RAND_1141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_733_im = _RAND_1142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_734_re = _RAND_1143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_734_im = _RAND_1144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_735_re = _RAND_1145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_735_im = _RAND_1146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_736_re = _RAND_1147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_736_im = _RAND_1148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_737_re = _RAND_1149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_737_im = _RAND_1150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_738_re = _RAND_1151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_738_im = _RAND_1152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_739_re = _RAND_1153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_739_im = _RAND_1154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_740_re = _RAND_1155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_740_im = _RAND_1156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_741_re = _RAND_1157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_741_im = _RAND_1158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_751_re = _RAND_1159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_751_im = _RAND_1160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_752_re = _RAND_1161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_752_im = _RAND_1162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_753_re = _RAND_1163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_753_im = _RAND_1164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_754_re = _RAND_1165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_754_im = _RAND_1166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_755_re = _RAND_1167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_755_im = _RAND_1168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_756_re = _RAND_1169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_756_im = _RAND_1170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_757_re = _RAND_1171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_757_im = _RAND_1172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_758_re = _RAND_1173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_758_im = _RAND_1174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_759_re = _RAND_1175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_759_im = _RAND_1176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_760_re = _RAND_1177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_760_im = _RAND_1178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_761_re = _RAND_1179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_761_im = _RAND_1180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_762_re = _RAND_1181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_762_im = _RAND_1182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_763_re = _RAND_1183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_763_im = _RAND_1184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_764_re = _RAND_1185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_764_im = _RAND_1186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_765_re = _RAND_1187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_765_im = _RAND_1188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_766_re = _RAND_1189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_766_im = _RAND_1190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_767_re = _RAND_1191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_767_im = _RAND_1192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_768_re = _RAND_1193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_768_im = _RAND_1194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_769_re = _RAND_1195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_769_im = _RAND_1196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_770_re = _RAND_1197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_770_im = _RAND_1198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_771_re = _RAND_1199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_771_im = _RAND_1200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_772_re = _RAND_1201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_772_im = _RAND_1202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_773_re = _RAND_1203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_773_im = _RAND_1204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_774_re = _RAND_1205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_774_im = _RAND_1206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_775_re = _RAND_1207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_775_im = _RAND_1208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_776_re = _RAND_1209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_776_im = _RAND_1210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_777_re = _RAND_1211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_777_im = _RAND_1212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_778_re = _RAND_1213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_778_im = _RAND_1214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_779_re = _RAND_1215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_779_im = _RAND_1216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_780_re = _RAND_1217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_780_im = _RAND_1218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_781_re = _RAND_1219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_781_im = _RAND_1220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_782_re = _RAND_1221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_782_im = _RAND_1222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_783_re = _RAND_1223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_783_im = _RAND_1224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_784_re = _RAND_1225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_784_im = _RAND_1226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_785_re = _RAND_1227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_785_im = _RAND_1228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_786_re = _RAND_1229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_786_im = _RAND_1230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_787_re = _RAND_1231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_787_im = _RAND_1232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_788_re = _RAND_1233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_788_im = _RAND_1234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_789_re = _RAND_1235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_789_im = _RAND_1236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_790_re = _RAND_1237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_790_im = _RAND_1238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_791_re = _RAND_1239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_791_im = _RAND_1240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_792_re = _RAND_1241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_792_im = _RAND_1242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_793_re = _RAND_1243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_793_im = _RAND_1244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_794_re = _RAND_1245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_794_im = _RAND_1246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_795_re = _RAND_1247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_795_im = _RAND_1248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_796_re = _RAND_1249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_796_im = _RAND_1250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_797_re = _RAND_1251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  _T_797_im = _RAND_1252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  _T_798_re = _RAND_1253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  _T_798_im = _RAND_1254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  _T_799_re = _RAND_1255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  _T_799_im = _RAND_1256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  _T_800_re = _RAND_1257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  _T_800_im = _RAND_1258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  _T_801_re = _RAND_1259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  _T_801_im = _RAND_1260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  _T_802_re = _RAND_1261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  _T_802_im = _RAND_1262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  _T_803_re = _RAND_1263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  _T_803_im = _RAND_1264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  _T_804_re = _RAND_1265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  _T_804_im = _RAND_1266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  _T_805_re = _RAND_1267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  _T_805_im = _RAND_1268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  _T_806_re = _RAND_1269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  _T_806_im = _RAND_1270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  _T_807_re = _RAND_1271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  _T_807_im = _RAND_1272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  _T_808_re = _RAND_1273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  _T_808_im = _RAND_1274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  _T_809_re = _RAND_1275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  _T_809_im = _RAND_1276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  _T_810_re = _RAND_1277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  _T_810_im = _RAND_1278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  _T_811_re = _RAND_1279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  _T_811_im = _RAND_1280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  _T_812_re = _RAND_1281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  _T_812_im = _RAND_1282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  _T_813_re = _RAND_1283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  _T_813_im = _RAND_1284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  _T_814_re = _RAND_1285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  _T_814_im = _RAND_1286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  _T_817_re = _RAND_1287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  _T_817_im = _RAND_1288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  _T_818_re = _RAND_1289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  _T_818_im = _RAND_1290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  _T_819_re = _RAND_1291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  _T_819_im = _RAND_1292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  _T_820_re = _RAND_1293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  _T_820_im = _RAND_1294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  _T_821_re = _RAND_1295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  _T_821_im = _RAND_1296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  _T_822_re = _RAND_1297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  _T_822_im = _RAND_1298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  _T_823_re = _RAND_1299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  _T_823_im = _RAND_1300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  _T_824_re = _RAND_1301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  _T_824_im = _RAND_1302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  _T_825_re = _RAND_1303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  _T_825_im = _RAND_1304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  _T_826_re = _RAND_1305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  _T_826_im = _RAND_1306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  _T_827_re = _RAND_1307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  _T_827_im = _RAND_1308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  _T_828_re = _RAND_1309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  _T_828_im = _RAND_1310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  _T_829_re = _RAND_1311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  _T_829_im = _RAND_1312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  _T_830_re = _RAND_1313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  _T_830_im = _RAND_1314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  _T_831_re = _RAND_1315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  _T_831_im = _RAND_1316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  _T_832_re = _RAND_1317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  _T_832_im = _RAND_1318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  _T_833_re = _RAND_1319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  _T_833_im = _RAND_1320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  _T_834_re = _RAND_1321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  _T_834_im = _RAND_1322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  _T_835_re = _RAND_1323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  _T_835_im = _RAND_1324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  _T_836_re = _RAND_1325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  _T_836_im = _RAND_1326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  _T_837_re = _RAND_1327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  _T_837_im = _RAND_1328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  _T_838_re = _RAND_1329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  _T_838_im = _RAND_1330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  _T_839_re = _RAND_1331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  _T_839_im = _RAND_1332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  _T_840_re = _RAND_1333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  _T_840_im = _RAND_1334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  _T_841_re = _RAND_1335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  _T_841_im = _RAND_1336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  _T_842_re = _RAND_1337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  _T_842_im = _RAND_1338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  _T_843_re = _RAND_1339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  _T_843_im = _RAND_1340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  _T_844_re = _RAND_1341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  _T_844_im = _RAND_1342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  _T_845_re = _RAND_1343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  _T_845_im = _RAND_1344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  _T_846_re = _RAND_1345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  _T_846_im = _RAND_1346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  _T_847_re = _RAND_1347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  _T_847_im = _RAND_1348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  _T_848_re = _RAND_1349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  _T_848_im = _RAND_1350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  _T_858_re = _RAND_1351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  _T_858_im = _RAND_1352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  _T_859_re = _RAND_1353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  _T_859_im = _RAND_1354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  _T_860_re = _RAND_1355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  _T_860_im = _RAND_1356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  _T_861_re = _RAND_1357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  _T_861_im = _RAND_1358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  _T_862_re = _RAND_1359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  _T_862_im = _RAND_1360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  _T_863_re = _RAND_1361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  _T_863_im = _RAND_1362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  _T_864_re = _RAND_1363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  _T_864_im = _RAND_1364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  _T_865_re = _RAND_1365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  _T_865_im = _RAND_1366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  _T_866_re = _RAND_1367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  _T_866_im = _RAND_1368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  _T_867_re = _RAND_1369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  _T_867_im = _RAND_1370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  _T_868_re = _RAND_1371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  _T_868_im = _RAND_1372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  _T_869_re = _RAND_1373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  _T_869_im = _RAND_1374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  _T_870_re = _RAND_1375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  _T_870_im = _RAND_1376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  _T_871_re = _RAND_1377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  _T_871_im = _RAND_1378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  _T_872_re = _RAND_1379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  _T_872_im = _RAND_1380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  _T_873_re = _RAND_1381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  _T_873_im = _RAND_1382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  _T_874_re = _RAND_1383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  _T_874_im = _RAND_1384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  _T_875_re = _RAND_1385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  _T_875_im = _RAND_1386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  _T_876_re = _RAND_1387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  _T_876_im = _RAND_1388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  _T_877_re = _RAND_1389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  _T_877_im = _RAND_1390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  _T_878_re = _RAND_1391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  _T_878_im = _RAND_1392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  _T_879_re = _RAND_1393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  _T_879_im = _RAND_1394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  _T_880_re = _RAND_1395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  _T_880_im = _RAND_1396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  _T_881_re = _RAND_1397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  _T_881_im = _RAND_1398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  _T_882_re = _RAND_1399[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  _T_882_im = _RAND_1400[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  _T_883_re = _RAND_1401[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  _T_883_im = _RAND_1402[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  _T_884_re = _RAND_1403[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  _T_884_im = _RAND_1404[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  _T_885_re = _RAND_1405[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  _T_885_im = _RAND_1406[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  _T_886_re = _RAND_1407[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  _T_886_im = _RAND_1408[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  _T_887_re = _RAND_1409[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  _T_887_im = _RAND_1410[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  _T_888_re = _RAND_1411[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  _T_888_im = _RAND_1412[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  _T_889_re = _RAND_1413[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  _T_889_im = _RAND_1414[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  _T_892_re = _RAND_1415[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  _T_892_im = _RAND_1416[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  _T_893_re = _RAND_1417[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  _T_893_im = _RAND_1418[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  _T_894_re = _RAND_1419[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  _T_894_im = _RAND_1420[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  _T_895_re = _RAND_1421[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  _T_895_im = _RAND_1422[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  _T_896_re = _RAND_1423[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  _T_896_im = _RAND_1424[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  _T_897_re = _RAND_1425[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  _T_897_im = _RAND_1426[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  _T_898_re = _RAND_1427[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  _T_898_im = _RAND_1428[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  _T_899_re = _RAND_1429[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  _T_899_im = _RAND_1430[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  _T_900_re = _RAND_1431[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  _T_900_im = _RAND_1432[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  _T_901_re = _RAND_1433[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  _T_901_im = _RAND_1434[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  _T_902_re = _RAND_1435[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  _T_902_im = _RAND_1436[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  _T_903_re = _RAND_1437[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  _T_903_im = _RAND_1438[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  _T_904_re = _RAND_1439[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  _T_904_im = _RAND_1440[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  _T_905_re = _RAND_1441[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  _T_905_im = _RAND_1442[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  _T_906_re = _RAND_1443[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  _T_906_im = _RAND_1444[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  _T_907_re = _RAND_1445[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  _T_907_im = _RAND_1446[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  _T_913_re = _RAND_1447[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  _T_913_im = _RAND_1448[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  _T_914_re = _RAND_1449[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  _T_914_im = _RAND_1450[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  _T_915_re = _RAND_1451[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  _T_915_im = _RAND_1452[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  _T_916_re = _RAND_1453[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  _T_916_im = _RAND_1454[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  _T_917_re = _RAND_1455[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  _T_917_im = _RAND_1456[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  _T_918_re = _RAND_1457[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  _T_918_im = _RAND_1458[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  _T_919_re = _RAND_1459[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  _T_919_im = _RAND_1460[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  _T_920_re = _RAND_1461[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  _T_920_im = _RAND_1462[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  _T_921_re = _RAND_1463[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  _T_921_im = _RAND_1464[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  _T_922_re = _RAND_1465[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  _T_922_im = _RAND_1466[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  _T_923_re = _RAND_1467[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  _T_923_im = _RAND_1468[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  _T_924_re = _RAND_1469[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  _T_924_im = _RAND_1470[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  _T_925_re = _RAND_1471[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  _T_925_im = _RAND_1472[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  _T_926_re = _RAND_1473[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  _T_926_im = _RAND_1474[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  _T_927_re = _RAND_1475[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  _T_927_im = _RAND_1476[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  _T_928_re = _RAND_1477[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  _T_928_im = _RAND_1478[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  _T_931_re = _RAND_1479[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  _T_931_im = _RAND_1480[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  _T_932_re = _RAND_1481[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  _T_932_im = _RAND_1482[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  _T_933_re = _RAND_1483[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  _T_933_im = _RAND_1484[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  _T_934_re = _RAND_1485[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  _T_934_im = _RAND_1486[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  _T_935_re = _RAND_1487[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  _T_935_im = _RAND_1488[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  _T_936_re = _RAND_1489[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  _T_936_im = _RAND_1490[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  _T_937_re = _RAND_1491[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  _T_937_im = _RAND_1492[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  _T_938_re = _RAND_1493[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  _T_938_im = _RAND_1494[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  _T_944_re = _RAND_1495[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  _T_944_im = _RAND_1496[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  _T_945_re = _RAND_1497[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  _T_945_im = _RAND_1498[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  _T_946_re = _RAND_1499[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  _T_946_im = _RAND_1500[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  _T_947_re = _RAND_1501[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  _T_947_im = _RAND_1502[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  _T_948_re = _RAND_1503[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  _T_948_im = _RAND_1504[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  _T_949_re = _RAND_1505[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  _T_949_im = _RAND_1506[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  _T_950_re = _RAND_1507[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  _T_950_im = _RAND_1508[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  _T_951_re = _RAND_1509[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  _T_951_im = _RAND_1510[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  _T_954_re = _RAND_1511[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  _T_954_im = _RAND_1512[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  _T_955_re = _RAND_1513[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  _T_955_im = _RAND_1514[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  _T_956_re = _RAND_1515[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  _T_956_im = _RAND_1516[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  _T_957_re = _RAND_1517[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  _T_957_im = _RAND_1518[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  _T_963_re = _RAND_1519[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  _T_963_im = _RAND_1520[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  _T_964_re = _RAND_1521[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  _T_964_im = _RAND_1522[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  _T_965_re = _RAND_1523[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  _T_965_im = _RAND_1524[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  _T_966_re = _RAND_1525[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  _T_966_im = _RAND_1526[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  _T_969_re = _RAND_1527[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  _T_969_im = _RAND_1528[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  _T_970_re = _RAND_1529[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  _T_970_im = _RAND_1530[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  _T_976_re = _RAND_1531[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  _T_976_im = _RAND_1532[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  _T_977_re = _RAND_1533[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  _T_977_im = _RAND_1534[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  _T_980_re = _RAND_1535[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  _T_980_im = _RAND_1536[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  out1D1_re = _RAND_1537[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  out1D1_im = _RAND_1538[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  _T_981_re = _RAND_1539[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  _T_981_im = _RAND_1540[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  _T_982_re = _RAND_1541[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  _T_982_im = _RAND_1542[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 9'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    cntD1 <= cnt;
    cntD2 <= cntD1;
    out1_0_re <= io_dIn_re;
    out1_0_im <= io_dIn_im;
    out2_0_re <= io_dIn_re;
    out2_0_im <= io_dIn_im;
    _T_153_re <= out1_0_re;
    _T_153_im <= out1_0_im;
    _T_154_re <= _T_153_re;
    _T_154_im <= _T_153_im;
    _T_155_re <= _T_154_re;
    _T_155_im <= _T_154_im;
    _T_156_re <= _T_155_re;
    _T_156_im <= _T_155_im;
    _T_157_re <= _T_156_re;
    _T_157_im <= _T_156_im;
    _T_158_re <= _T_157_re;
    _T_158_im <= _T_157_im;
    _T_159_re <= _T_158_re;
    _T_159_im <= _T_158_im;
    _T_160_re <= _T_159_re;
    _T_160_im <= _T_159_im;
    _T_161_re <= _T_160_re;
    _T_161_im <= _T_160_im;
    _T_162_re <= _T_161_re;
    _T_162_im <= _T_161_im;
    _T_163_re <= _T_162_re;
    _T_163_im <= _T_162_im;
    _T_164_re <= _T_163_re;
    _T_164_im <= _T_163_im;
    _T_165_re <= _T_164_re;
    _T_165_im <= _T_164_im;
    _T_166_re <= _T_165_re;
    _T_166_im <= _T_165_im;
    _T_167_re <= _T_166_re;
    _T_167_im <= _T_166_im;
    _T_168_re <= _T_167_re;
    _T_168_im <= _T_167_im;
    _T_169_re <= _T_168_re;
    _T_169_im <= _T_168_im;
    _T_170_re <= _T_169_re;
    _T_170_im <= _T_169_im;
    _T_171_re <= _T_170_re;
    _T_171_im <= _T_170_im;
    _T_172_re <= _T_171_re;
    _T_172_im <= _T_171_im;
    _T_173_re <= _T_172_re;
    _T_173_im <= _T_172_im;
    _T_174_re <= _T_173_re;
    _T_174_im <= _T_173_im;
    _T_175_re <= _T_174_re;
    _T_175_im <= _T_174_im;
    _T_176_re <= _T_175_re;
    _T_176_im <= _T_175_im;
    _T_177_re <= _T_176_re;
    _T_177_im <= _T_176_im;
    _T_178_re <= _T_177_re;
    _T_178_im <= _T_177_im;
    _T_179_re <= _T_178_re;
    _T_179_im <= _T_178_im;
    _T_180_re <= _T_179_re;
    _T_180_im <= _T_179_im;
    _T_181_re <= _T_180_re;
    _T_181_im <= _T_180_im;
    _T_182_re <= _T_181_re;
    _T_182_im <= _T_181_im;
    _T_183_re <= _T_182_re;
    _T_183_im <= _T_182_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_325_re <= _T_324_re;
    _T_325_im <= _T_324_im;
    _T_326_re <= _T_325_re;
    _T_326_im <= _T_325_im;
    _T_327_re <= _T_326_re;
    _T_327_im <= _T_326_im;
    _T_328_re <= _T_327_re;
    _T_328_im <= _T_327_im;
    _T_329_re <= _T_328_re;
    _T_329_im <= _T_328_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_393_re <= _T_392_re;
    _T_393_im <= _T_392_im;
    _T_394_re <= _T_393_re;
    _T_394_im <= _T_393_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_402_re <= _T_401_re;
    _T_402_im <= _T_401_im;
    _T_403_re <= _T_402_re;
    _T_403_im <= _T_402_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_406_re <= _T_405_re;
    _T_406_im <= _T_405_im;
    _T_407_re <= _T_406_re;
    _T_407_im <= _T_406_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_411_re <= Butterfly_io_out2_re;
    _T_411_im <= Butterfly_io_out2_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_533_re <= _T_532_re;
    _T_533_im <= _T_532_im;
    _T_534_re <= _T_533_re;
    _T_534_im <= _T_533_im;
    _T_535_re <= _T_534_re;
    _T_535_im <= _T_534_im;
    _T_536_re <= _T_535_re;
    _T_536_im <= _T_535_im;
    _T_537_re <= _T_536_re;
    _T_537_im <= _T_536_im;
    _T_538_re <= _T_537_re;
    _T_538_im <= _T_537_im;
    _T_548_re <= Switch_io_out1_re;
    _T_548_im <= Switch_io_out1_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_663_re <= _T_662_re;
    _T_663_im <= _T_662_im;
    _T_664_re <= _T_663_re;
    _T_664_im <= _T_663_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_671_re <= _T_670_re;
    _T_671_im <= _T_670_im;
    _T_672_re <= _T_671_re;
    _T_672_im <= _T_671_im;
    _T_673_re <= _T_672_re;
    _T_673_im <= _T_672_im;
    _T_674_re <= _T_673_re;
    _T_674_im <= _T_673_im;
    _T_675_re <= _T_674_re;
    _T_675_im <= _T_674_im;
    _T_678_re <= Butterfly_1_io_out2_re;
    _T_678_im <= Butterfly_1_io_out2_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_728_re <= _T_727_re;
    _T_728_im <= _T_727_im;
    _T_729_re <= _T_728_re;
    _T_729_im <= _T_728_im;
    _T_730_re <= _T_729_re;
    _T_730_im <= _T_729_im;
    _T_731_re <= _T_730_re;
    _T_731_im <= _T_730_im;
    _T_732_re <= _T_731_re;
    _T_732_im <= _T_731_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_736_re <= _T_735_re;
    _T_736_im <= _T_735_im;
    _T_737_re <= _T_736_re;
    _T_737_im <= _T_736_im;
    _T_738_re <= _T_737_re;
    _T_738_im <= _T_737_im;
    _T_739_re <= _T_738_re;
    _T_739_im <= _T_738_im;
    _T_740_re <= _T_739_re;
    _T_740_im <= _T_739_im;
    _T_741_re <= _T_740_re;
    _T_741_im <= _T_740_im;
    _T_751_re <= Switch_1_io_out1_re;
    _T_751_im <= Switch_1_io_out1_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_796_re <= _T_795_re;
    _T_796_im <= _T_795_im;
    _T_797_re <= _T_796_re;
    _T_797_im <= _T_796_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_808_re <= _T_807_re;
    _T_808_im <= _T_807_im;
    _T_809_re <= _T_808_re;
    _T_809_im <= _T_808_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_811_re <= _T_810_re;
    _T_811_im <= _T_810_im;
    _T_812_re <= _T_811_re;
    _T_812_im <= _T_811_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_817_re <= Butterfly_2_io_out2_re;
    _T_817_im <= Butterfly_2_io_out2_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_829_re <= _T_828_re;
    _T_829_im <= _T_828_im;
    _T_830_re <= _T_829_re;
    _T_830_im <= _T_829_im;
    _T_831_re <= _T_830_re;
    _T_831_im <= _T_830_im;
    _T_832_re <= _T_831_re;
    _T_832_im <= _T_831_im;
    _T_833_re <= _T_832_re;
    _T_833_im <= _T_832_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_841_re <= _T_840_re;
    _T_841_im <= _T_840_im;
    _T_842_re <= _T_841_re;
    _T_842_im <= _T_841_im;
    _T_843_re <= _T_842_re;
    _T_843_im <= _T_842_im;
    _T_844_re <= _T_843_re;
    _T_844_im <= _T_843_im;
    _T_845_re <= _T_844_re;
    _T_845_im <= _T_844_im;
    _T_846_re <= _T_845_re;
    _T_846_im <= _T_845_im;
    _T_847_re <= _T_846_re;
    _T_847_im <= _T_846_im;
    _T_848_re <= _T_847_re;
    _T_848_im <= _T_847_im;
    _T_858_re <= Switch_2_io_out1_re;
    _T_858_im <= Switch_2_io_out1_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_865_re <= _T_864_re;
    _T_865_im <= _T_864_im;
    _T_866_re <= _T_865_re;
    _T_866_im <= _T_865_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_881_re <= _T_880_re;
    _T_881_im <= _T_880_im;
    _T_882_re <= _T_881_re;
    _T_882_im <= _T_881_im;
    _T_883_re <= _T_882_re;
    _T_883_im <= _T_882_im;
    _T_884_re <= _T_883_re;
    _T_884_im <= _T_883_im;
    _T_885_re <= _T_884_re;
    _T_885_im <= _T_884_im;
    _T_886_re <= _T_885_re;
    _T_886_im <= _T_885_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_892_re <= Butterfly_3_io_out2_re;
    _T_892_im <= Butterfly_3_io_out2_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_898_re <= _T_897_re;
    _T_898_im <= _T_897_im;
    _T_899_re <= _T_898_re;
    _T_899_im <= _T_898_im;
    _T_900_re <= _T_899_re;
    _T_900_im <= _T_899_im;
    _T_901_re <= _T_900_re;
    _T_901_im <= _T_900_im;
    _T_902_re <= _T_901_re;
    _T_902_im <= _T_901_im;
    _T_903_re <= _T_902_re;
    _T_903_im <= _T_902_im;
    _T_904_re <= _T_903_re;
    _T_904_im <= _T_903_im;
    _T_905_re <= _T_904_re;
    _T_905_im <= _T_904_im;
    _T_906_re <= _T_905_re;
    _T_906_im <= _T_905_im;
    _T_907_re <= _T_906_re;
    _T_907_im <= _T_906_im;
    _T_913_re <= Switch_3_io_out1_re;
    _T_913_im <= Switch_3_io_out1_im;
    _T_914_re <= _T_913_re;
    _T_914_im <= _T_913_im;
    _T_915_re <= _T_914_re;
    _T_915_im <= _T_914_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_922_re <= _T_921_re;
    _T_922_im <= _T_921_im;
    _T_923_re <= _T_922_re;
    _T_923_im <= _T_922_im;
    _T_924_re <= _T_923_re;
    _T_924_im <= _T_923_im;
    _T_925_re <= _T_924_re;
    _T_925_im <= _T_924_im;
    _T_926_re <= _T_925_re;
    _T_926_im <= _T_925_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_928_re <= _T_927_re;
    _T_928_im <= _T_927_im;
    _T_931_re <= Butterfly_4_io_out2_re;
    _T_931_im <= Butterfly_4_io_out2_im;
    _T_932_re <= _T_931_re;
    _T_932_im <= _T_931_im;
    _T_933_re <= _T_932_re;
    _T_933_im <= _T_932_im;
    _T_934_re <= _T_933_re;
    _T_934_im <= _T_933_im;
    _T_935_re <= _T_934_re;
    _T_935_im <= _T_934_im;
    _T_936_re <= _T_935_re;
    _T_936_im <= _T_935_im;
    _T_937_re <= _T_936_re;
    _T_937_im <= _T_936_im;
    _T_938_re <= _T_937_re;
    _T_938_im <= _T_937_im;
    _T_944_re <= Switch_4_io_out1_re;
    _T_944_im <= Switch_4_io_out1_im;
    _T_945_re <= _T_944_re;
    _T_945_im <= _T_944_im;
    _T_946_re <= _T_945_re;
    _T_946_im <= _T_945_im;
    _T_947_re <= _T_946_re;
    _T_947_im <= _T_946_im;
    _T_948_re <= _T_947_re;
    _T_948_im <= _T_947_im;
    _T_949_re <= _T_948_re;
    _T_949_im <= _T_948_im;
    _T_950_re <= _T_949_re;
    _T_950_im <= _T_949_im;
    _T_951_re <= _T_950_re;
    _T_951_im <= _T_950_im;
    _T_954_re <= Butterfly_5_io_out2_re;
    _T_954_im <= Butterfly_5_io_out2_im;
    _T_955_re <= _T_954_re;
    _T_955_im <= _T_954_im;
    _T_956_re <= _T_955_re;
    _T_956_im <= _T_955_im;
    _T_957_re <= _T_956_re;
    _T_957_im <= _T_956_im;
    _T_963_re <= Switch_5_io_out1_re;
    _T_963_im <= Switch_5_io_out1_im;
    _T_964_re <= _T_963_re;
    _T_964_im <= _T_963_im;
    _T_965_re <= _T_964_re;
    _T_965_im <= _T_964_im;
    _T_966_re <= _T_965_re;
    _T_966_im <= _T_965_im;
    _T_969_re <= Butterfly_6_io_out2_re;
    _T_969_im <= Butterfly_6_io_out2_im;
    _T_970_re <= _T_969_re;
    _T_970_im <= _T_969_im;
    _T_976_re <= Switch_6_io_out1_re;
    _T_976_im <= Switch_6_io_out1_im;
    _T_977_re <= _T_976_re;
    _T_977_im <= _T_976_im;
    _T_980_re <= Butterfly_7_io_out2_re;
    _T_980_im <= Butterfly_7_io_out2_im;
    out1D1_re <= Switch_7_io_out1_re;
    out1D1_im <= Switch_7_io_out1_im;
    _T_981_re <= ComplexAdd_io_res_re;
    _T_981_im <= ComplexAdd_io_res_im;
    _T_982_re <= ComplexSub_io_res_re;
    _T_982_im <= ComplexSub_io_res_im;
  end
endmodule
